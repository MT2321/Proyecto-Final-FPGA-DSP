LIBRARY ieee;
USE ieee.STD_LOGIC_1164.ALL;
USE ieee.std_logic_unsigned.all;
USE ieee.numeric_std.ALL;

ENTITY LUT IS
	PORT(
		table_in:	IN STD_LOGIC_VECTOR(11 DOWNTO 0);
		table_out:	OUT INTEGER RANGE 0 TO 4095
	);
END LUT;

ARCHITECTURE Behavior OF LUT IS
BEGIN

	PROCESS(table_in)
	BEGIN
		CASE table_in IS
			WHEN "000000000000" => table_out <= 0;
			WHEN "000000000001" => table_out <= 1;
			WHEN "000000000010" => table_out <= 342;
			WHEN "000000000011" => table_out <= 541;
			WHEN "000000000100" => table_out <= 683;
			WHEN "000000000101" => table_out <= 793;
			WHEN "000000000110" => table_out <= 882;
			WHEN "000000000111" => table_out <= 958;
			WHEN "000000001000" => table_out <= 1024;
			WHEN "000000001001" => table_out <= 1082;
			WHEN "000000001010" => table_out <= 1134;
			WHEN "000000001011" => table_out <= 1181;
			WHEN "000000001100" => table_out <= 1224;
			WHEN "000000001101" => table_out <= 1263;
			WHEN "000000001110" => table_out <= 1299;
			WHEN "000000001111" => table_out <= 1333;
			WHEN "000000010000" => table_out <= 1365;
			WHEN "000000010001" => table_out <= 1395;
			WHEN "000000010010" => table_out <= 1423;
			WHEN "000000010011" => table_out <= 1450;
			WHEN "000000010100" => table_out <= 1475;
			WHEN "000000010101" => table_out <= 1499;
			WHEN "000000010110" => table_out <= 1522;
			WHEN "000000010111" => table_out <= 1544;
			WHEN "000000011000" => table_out <= 1565;
			WHEN "000000011001" => table_out <= 1585;
			WHEN "000000011010" => table_out <= 1604;
			WHEN "000000011011" => table_out <= 1623;
			WHEN "000000011100" => table_out <= 1641;
			WHEN "000000011101" => table_out <= 1658;
			WHEN "000000011110" => table_out <= 1675;
			WHEN "000000011111" => table_out <= 1691;
			WHEN "000000100000" => table_out <= 1706;
			WHEN "000000100001" => table_out <= 1722;
			WHEN "000000100010" => table_out <= 1736;
			WHEN "000000100011" => table_out <= 1750;
			WHEN "000000100100" => table_out <= 1764;
			WHEN "000000100101" => table_out <= 1778;
			WHEN "000000100110" => table_out <= 1791;
			WHEN "000000100111" => table_out <= 1804;
			WHEN "000000101000" => table_out <= 1816;
			WHEN "000000101001" => table_out <= 1828;
			WHEN "000000101010" => table_out <= 1840;
			WHEN "000000101011" => table_out <= 1852;
			WHEN "000000101100" => table_out <= 1863;
			WHEN "000000101101" => table_out <= 1874;
			WHEN "000000101110" => table_out <= 1885;
			WHEN "000000101111" => table_out <= 1896;
			WHEN "000000110000" => table_out <= 1906;
			WHEN "000000110001" => table_out <= 1916;
			WHEN "000000110010" => table_out <= 1926;
			WHEN "000000110011" => table_out <= 1936;
			WHEN "000000110100" => table_out <= 1945;
			WHEN "000000110101" => table_out <= 1955;
			WHEN "000000110110" => table_out <= 1964;
			WHEN "000000110111" => table_out <= 1973;
			WHEN "000000111000" => table_out <= 1982;
			WHEN "000000111001" => table_out <= 1991;
			WHEN "000000111010" => table_out <= 1999;
			WHEN "000000111011" => table_out <= 2008;
			WHEN "000000111100" => table_out <= 2016;
			WHEN "000000111101" => table_out <= 2024;
			WHEN "000000111110" => table_out <= 2032;
			WHEN "000000111111" => table_out <= 2040;
			WHEN "000001000000" => table_out <= 2048;
			WHEN "000001000001" => table_out <= 2055;
			WHEN "000001000010" => table_out <= 2063;
			WHEN "000001000011" => table_out <= 2070;
			WHEN "000001000100" => table_out <= 2077;
			WHEN "000001000101" => table_out <= 2085;
			WHEN "000001000110" => table_out <= 2092;
			WHEN "000001000111" => table_out <= 2099;
			WHEN "000001001000" => table_out <= 2106;
			WHEN "000001001001" => table_out <= 2112;
			WHEN "000001001010" => table_out <= 2119;
			WHEN "000001001011" => table_out <= 2126;
			WHEN "000001001100" => table_out <= 2132;
			WHEN "000001001101" => table_out <= 2139;
			WHEN "000001001110" => table_out <= 2145;
			WHEN "000001001111" => table_out <= 2151;
			WHEN "000001010000" => table_out <= 2157;
			WHEN "000001010001" => table_out <= 2164;
			WHEN "000001010010" => table_out <= 2170;
			WHEN "000001010011" => table_out <= 2176;
			WHEN "000001010100" => table_out <= 2181;
			WHEN "000001010101" => table_out <= 2187;
			WHEN "000001010110" => table_out <= 2193;
			WHEN "000001010111" => table_out <= 2199;
			WHEN "000001011000" => table_out <= 2204;
			WHEN "000001011001" => table_out <= 2210;
			WHEN "000001011010" => table_out <= 2215;
			WHEN "000001011011" => table_out <= 2221;
			WHEN "000001011100" => table_out <= 2226;
			WHEN "000001011101" => table_out <= 2232;
			WHEN "000001011110" => table_out <= 2237;
			WHEN "000001011111" => table_out <= 2242;
			WHEN "000001100000" => table_out <= 2247;
			WHEN "000001100001" => table_out <= 2252;
			WHEN "000001100010" => table_out <= 2257;
			WHEN "000001100011" => table_out <= 2262;
			WHEN "000001100100" => table_out <= 2267;
			WHEN "000001100101" => table_out <= 2272;
			WHEN "000001100110" => table_out <= 2277;
			WHEN "000001100111" => table_out <= 2282;
			WHEN "000001101000" => table_out <= 2287;
			WHEN "000001101001" => table_out <= 2291;
			WHEN "000001101010" => table_out <= 2296;
			WHEN "000001101011" => table_out <= 2301;
			WHEN "000001101100" => table_out <= 2305;
			WHEN "000001101101" => table_out <= 2310;
			WHEN "000001101110" => table_out <= 2314;
			WHEN "000001101111" => table_out <= 2319;
			WHEN "000001110000" => table_out <= 2323;
			WHEN "000001110001" => table_out <= 2327;
			WHEN "000001110010" => table_out <= 2332;
			WHEN "000001110011" => table_out <= 2336;
			WHEN "000001110100" => table_out <= 2340;
			WHEN "000001110101" => table_out <= 2345;
			WHEN "000001110110" => table_out <= 2349;
			WHEN "000001110111" => table_out <= 2353;
			WHEN "000001111000" => table_out <= 2357;
			WHEN "000001111001" => table_out <= 2361;
			WHEN "000001111010" => table_out <= 2365;
			WHEN "000001111011" => table_out <= 2369;
			WHEN "000001111100" => table_out <= 2373;
			WHEN "000001111101" => table_out <= 2377;
			WHEN "000001111110" => table_out <= 2381;
			WHEN "000001111111" => table_out <= 2385;
			WHEN "000010000000" => table_out <= 2389;
			WHEN "000010000001" => table_out <= 2393;
			WHEN "000010000010" => table_out <= 2396;
			WHEN "000010000011" => table_out <= 2400;
			WHEN "000010000100" => table_out <= 2404;
			WHEN "000010000101" => table_out <= 2408;
			WHEN "000010000110" => table_out <= 2411;
			WHEN "000010000111" => table_out <= 2415;
			WHEN "000010001000" => table_out <= 2419;
			WHEN "000010001001" => table_out <= 2422;
			WHEN "000010001010" => table_out <= 2426;
			WHEN "000010001011" => table_out <= 2429;
			WHEN "000010001100" => table_out <= 2433;
			WHEN "000010001101" => table_out <= 2436;
			WHEN "000010001110" => table_out <= 2440;
			WHEN "000010001111" => table_out <= 2443;
			WHEN "000010010000" => table_out <= 2447;
			WHEN "000010010001" => table_out <= 2450;
			WHEN "000010010010" => table_out <= 2454;
			WHEN "000010010011" => table_out <= 2457;
			WHEN "000010010100" => table_out <= 2460;
			WHEN "000010010101" => table_out <= 2464;
			WHEN "000010010110" => table_out <= 2467;
			WHEN "000010010111" => table_out <= 2470;
			WHEN "000010011000" => table_out <= 2473;
			WHEN "000010011001" => table_out <= 2477;
			WHEN "000010011010" => table_out <= 2480;
			WHEN "000010011011" => table_out <= 2483;
			WHEN "000010011100" => table_out <= 2486;
			WHEN "000010011101" => table_out <= 2489;
			WHEN "000010011110" => table_out <= 2492;
			WHEN "000010011111" => table_out <= 2495;
			WHEN "000010100000" => table_out <= 2499;
			WHEN "000010100001" => table_out <= 2502;
			WHEN "000010100010" => table_out <= 2505;
			WHEN "000010100011" => table_out <= 2508;
			WHEN "000010100100" => table_out <= 2511;
			WHEN "000010100101" => table_out <= 2514;
			WHEN "000010100110" => table_out <= 2517;
			WHEN "000010100111" => table_out <= 2520;
			WHEN "000010101000" => table_out <= 2523;
			WHEN "000010101001" => table_out <= 2526;
			WHEN "000010101010" => table_out <= 2528;
			WHEN "000010101011" => table_out <= 2531;
			WHEN "000010101100" => table_out <= 2534;
			WHEN "000010101101" => table_out <= 2537;
			WHEN "000010101110" => table_out <= 2540;
			WHEN "000010101111" => table_out <= 2543;
			WHEN "000010110000" => table_out <= 2545;
			WHEN "000010110001" => table_out <= 2548;
			WHEN "000010110010" => table_out <= 2551;
			WHEN "000010110011" => table_out <= 2554;
			WHEN "000010110100" => table_out <= 2557;
			WHEN "000010110101" => table_out <= 2559;
			WHEN "000010110110" => table_out <= 2562;
			WHEN "000010110111" => table_out <= 2565;
			WHEN "000010111000" => table_out <= 2567;
			WHEN "000010111001" => table_out <= 2570;
			WHEN "000010111010" => table_out <= 2573;
			WHEN "000010111011" => table_out <= 2575;
			WHEN "000010111100" => table_out <= 2578;
			WHEN "000010111101" => table_out <= 2581;
			WHEN "000010111110" => table_out <= 2583;
			WHEN "000010111111" => table_out <= 2586;
			WHEN "000011000000" => table_out <= 2588;
			WHEN "000011000001" => table_out <= 2591;
			WHEN "000011000010" => table_out <= 2593;
			WHEN "000011000011" => table_out <= 2596;
			WHEN "000011000100" => table_out <= 2598;
			WHEN "000011000101" => table_out <= 2601;
			WHEN "000011000110" => table_out <= 2603;
			WHEN "000011000111" => table_out <= 2606;
			WHEN "000011001000" => table_out <= 2608;
			WHEN "000011001001" => table_out <= 2611;
			WHEN "000011001010" => table_out <= 2613;
			WHEN "000011001011" => table_out <= 2616;
			WHEN "000011001100" => table_out <= 2618;
			WHEN "000011001101" => table_out <= 2621;
			WHEN "000011001110" => table_out <= 2623;
			WHEN "000011001111" => table_out <= 2625;
			WHEN "000011010000" => table_out <= 2628;
			WHEN "000011010001" => table_out <= 2630;
			WHEN "000011010010" => table_out <= 2632;
			WHEN "000011010011" => table_out <= 2635;
			WHEN "000011010100" => table_out <= 2637;
			WHEN "000011010101" => table_out <= 2639;
			WHEN "000011010110" => table_out <= 2642;
			WHEN "000011010111" => table_out <= 2644;
			WHEN "000011011000" => table_out <= 2646;
			WHEN "000011011001" => table_out <= 2649;
			WHEN "000011011010" => table_out <= 2651;
			WHEN "000011011011" => table_out <= 2653;
			WHEN "000011011100" => table_out <= 2655;
			WHEN "000011011101" => table_out <= 2658;
			WHEN "000011011110" => table_out <= 2660;
			WHEN "000011011111" => table_out <= 2662;
			WHEN "000011100000" => table_out <= 2664;
			WHEN "000011100001" => table_out <= 2666;
			WHEN "000011100010" => table_out <= 2669;
			WHEN "000011100011" => table_out <= 2671;
			WHEN "000011100100" => table_out <= 2673;
			WHEN "000011100101" => table_out <= 2675;
			WHEN "000011100110" => table_out <= 2677;
			WHEN "000011100111" => table_out <= 2679;
			WHEN "000011101000" => table_out <= 2681;
			WHEN "000011101001" => table_out <= 2684;
			WHEN "000011101010" => table_out <= 2686;
			WHEN "000011101011" => table_out <= 2688;
			WHEN "000011101100" => table_out <= 2690;
			WHEN "000011101101" => table_out <= 2692;
			WHEN "000011101110" => table_out <= 2694;
			WHEN "000011101111" => table_out <= 2696;
			WHEN "000011110000" => table_out <= 2698;
			WHEN "000011110001" => table_out <= 2700;
			WHEN "000011110010" => table_out <= 2702;
			WHEN "000011110011" => table_out <= 2704;
			WHEN "000011110100" => table_out <= 2706;
			WHEN "000011110101" => table_out <= 2708;
			WHEN "000011110110" => table_out <= 2710;
			WHEN "000011110111" => table_out <= 2712;
			WHEN "000011111000" => table_out <= 2714;
			WHEN "000011111001" => table_out <= 2716;
			WHEN "000011111010" => table_out <= 2718;
			WHEN "000011111011" => table_out <= 2720;
			WHEN "000011111100" => table_out <= 2722;
			WHEN "000011111101" => table_out <= 2724;
			WHEN "000011111110" => table_out <= 2726;
			WHEN "000011111111" => table_out <= 2728;
			WHEN "000100000000" => table_out <= 2730;
			WHEN "000100000001" => table_out <= 2732;
			WHEN "000100000010" => table_out <= 2734;
			WHEN "000100000011" => table_out <= 2736;
			WHEN "000100000100" => table_out <= 2738;
			WHEN "000100000101" => table_out <= 2739;
			WHEN "000100000110" => table_out <= 2741;
			WHEN "000100000111" => table_out <= 2743;
			WHEN "000100001000" => table_out <= 2745;
			WHEN "000100001001" => table_out <= 2747;
			WHEN "000100001010" => table_out <= 2749;
			WHEN "000100001011" => table_out <= 2751;
			WHEN "000100001100" => table_out <= 2752;
			WHEN "000100001101" => table_out <= 2754;
			WHEN "000100001110" => table_out <= 2756;
			WHEN "000100001111" => table_out <= 2758;
			WHEN "000100010000" => table_out <= 2760;
			WHEN "000100010001" => table_out <= 2762;
			WHEN "000100010010" => table_out <= 2763;
			WHEN "000100010011" => table_out <= 2765;
			WHEN "000100010100" => table_out <= 2767;
			WHEN "000100010101" => table_out <= 2769;
			WHEN "000100010110" => table_out <= 2770;
			WHEN "000100010111" => table_out <= 2772;
			WHEN "000100011000" => table_out <= 2774;
			WHEN "000100011001" => table_out <= 2776;
			WHEN "000100011010" => table_out <= 2778;
			WHEN "000100011011" => table_out <= 2779;
			WHEN "000100011100" => table_out <= 2781;
			WHEN "000100011101" => table_out <= 2783;
			WHEN "000100011110" => table_out <= 2784;
			WHEN "000100011111" => table_out <= 2786;
			WHEN "000100100000" => table_out <= 2788;
			WHEN "000100100001" => table_out <= 2790;
			WHEN "000100100010" => table_out <= 2791;
			WHEN "000100100011" => table_out <= 2793;
			WHEN "000100100100" => table_out <= 2795;
			WHEN "000100100101" => table_out <= 2796;
			WHEN "000100100110" => table_out <= 2798;
			WHEN "000100100111" => table_out <= 2800;
			WHEN "000100101000" => table_out <= 2801;
			WHEN "000100101001" => table_out <= 2803;
			WHEN "000100101010" => table_out <= 2805;
			WHEN "000100101011" => table_out <= 2806;
			WHEN "000100101100" => table_out <= 2808;
			WHEN "000100101101" => table_out <= 2810;
			WHEN "000100101110" => table_out <= 2811;
			WHEN "000100101111" => table_out <= 2813;
			WHEN "000100110000" => table_out <= 2815;
			WHEN "000100110001" => table_out <= 2816;
			WHEN "000100110010" => table_out <= 2818;
			WHEN "000100110011" => table_out <= 2819;
			WHEN "000100110100" => table_out <= 2821;
			WHEN "000100110101" => table_out <= 2823;
			WHEN "000100110110" => table_out <= 2824;
			WHEN "000100110111" => table_out <= 2826;
			WHEN "000100111000" => table_out <= 2827;
			WHEN "000100111001" => table_out <= 2829;
			WHEN "000100111010" => table_out <= 2830;
			WHEN "000100111011" => table_out <= 2832;
			WHEN "000100111100" => table_out <= 2834;
			WHEN "000100111101" => table_out <= 2835;
			WHEN "000100111110" => table_out <= 2837;
			WHEN "000100111111" => table_out <= 2838;
			WHEN "000101000000" => table_out <= 2840;
			WHEN "000101000001" => table_out <= 2841;
			WHEN "000101000010" => table_out <= 2843;
			WHEN "000101000011" => table_out <= 2844;
			WHEN "000101000100" => table_out <= 2846;
			WHEN "000101000101" => table_out <= 2847;
			WHEN "000101000110" => table_out <= 2849;
			WHEN "000101000111" => table_out <= 2850;
			WHEN "000101001000" => table_out <= 2852;
			WHEN "000101001001" => table_out <= 2853;
			WHEN "000101001010" => table_out <= 2855;
			WHEN "000101001011" => table_out <= 2856;
			WHEN "000101001100" => table_out <= 2858;
			WHEN "000101001101" => table_out <= 2859;
			WHEN "000101001110" => table_out <= 2861;
			WHEN "000101001111" => table_out <= 2862;
			WHEN "000101010000" => table_out <= 2864;
			WHEN "000101010001" => table_out <= 2865;
			WHEN "000101010010" => table_out <= 2867;
			WHEN "000101010011" => table_out <= 2868;
			WHEN "000101010100" => table_out <= 2870;
			WHEN "000101010101" => table_out <= 2871;
			WHEN "000101010110" => table_out <= 2872;
			WHEN "000101010111" => table_out <= 2874;
			WHEN "000101011000" => table_out <= 2875;
			WHEN "000101011001" => table_out <= 2877;
			WHEN "000101011010" => table_out <= 2878;
			WHEN "000101011011" => table_out <= 2880;
			WHEN "000101011100" => table_out <= 2881;
			WHEN "000101011101" => table_out <= 2882;
			WHEN "000101011110" => table_out <= 2884;
			WHEN "000101011111" => table_out <= 2885;
			WHEN "000101100000" => table_out <= 2887;
			WHEN "000101100001" => table_out <= 2888;
			WHEN "000101100010" => table_out <= 2889;
			WHEN "000101100011" => table_out <= 2891;
			WHEN "000101100100" => table_out <= 2892;
			WHEN "000101100101" => table_out <= 2894;
			WHEN "000101100110" => table_out <= 2895;
			WHEN "000101100111" => table_out <= 2896;
			WHEN "000101101000" => table_out <= 2898;
			WHEN "000101101001" => table_out <= 2899;
			WHEN "000101101010" => table_out <= 2900;
			WHEN "000101101011" => table_out <= 2902;
			WHEN "000101101100" => table_out <= 2903;
			WHEN "000101101101" => table_out <= 2905;
			WHEN "000101101110" => table_out <= 2906;
			WHEN "000101101111" => table_out <= 2907;
			WHEN "000101110000" => table_out <= 2909;
			WHEN "000101110001" => table_out <= 2910;
			WHEN "000101110010" => table_out <= 2911;
			WHEN "000101110011" => table_out <= 2913;
			WHEN "000101110100" => table_out <= 2914;
			WHEN "000101110101" => table_out <= 2915;
			WHEN "000101110110" => table_out <= 2917;
			WHEN "000101110111" => table_out <= 2918;
			WHEN "000101111000" => table_out <= 2919;
			WHEN "000101111001" => table_out <= 2920;
			WHEN "000101111010" => table_out <= 2922;
			WHEN "000101111011" => table_out <= 2923;
			WHEN "000101111100" => table_out <= 2924;
			WHEN "000101111101" => table_out <= 2926;
			WHEN "000101111110" => table_out <= 2927;
			WHEN "000101111111" => table_out <= 2928;
			WHEN "000110000000" => table_out <= 2929;
			WHEN "000110000001" => table_out <= 2931;
			WHEN "000110000010" => table_out <= 2932;
			WHEN "000110000011" => table_out <= 2933;
			WHEN "000110000100" => table_out <= 2935;
			WHEN "000110000101" => table_out <= 2936;
			WHEN "000110000110" => table_out <= 2937;
			WHEN "000110000111" => table_out <= 2938;
			WHEN "000110001000" => table_out <= 2940;
			WHEN "000110001001" => table_out <= 2941;
			WHEN "000110001010" => table_out <= 2942;
			WHEN "000110001011" => table_out <= 2943;
			WHEN "000110001100" => table_out <= 2945;
			WHEN "000110001101" => table_out <= 2946;
			WHEN "000110001110" => table_out <= 2947;
			WHEN "000110001111" => table_out <= 2948;
			WHEN "000110010000" => table_out <= 2950;
			WHEN "000110010001" => table_out <= 2951;
			WHEN "000110010010" => table_out <= 2952;
			WHEN "000110010011" => table_out <= 2953;
			WHEN "000110010100" => table_out <= 2954;
			WHEN "000110010101" => table_out <= 2956;
			WHEN "000110010110" => table_out <= 2957;
			WHEN "000110010111" => table_out <= 2958;
			WHEN "000110011000" => table_out <= 2959;
			WHEN "000110011001" => table_out <= 2961;
			WHEN "000110011010" => table_out <= 2962;
			WHEN "000110011011" => table_out <= 2963;
			WHEN "000110011100" => table_out <= 2964;
			WHEN "000110011101" => table_out <= 2965;
			WHEN "000110011110" => table_out <= 2967;
			WHEN "000110011111" => table_out <= 2968;
			WHEN "000110100000" => table_out <= 2969;
			WHEN "000110100001" => table_out <= 2970;
			WHEN "000110100010" => table_out <= 2971;
			WHEN "000110100011" => table_out <= 2972;
			WHEN "000110100100" => table_out <= 2974;
			WHEN "000110100101" => table_out <= 2975;
			WHEN "000110100110" => table_out <= 2976;
			WHEN "000110100111" => table_out <= 2977;
			WHEN "000110101000" => table_out <= 2978;
			WHEN "000110101001" => table_out <= 2979;
			WHEN "000110101010" => table_out <= 2981;
			WHEN "000110101011" => table_out <= 2982;
			WHEN "000110101100" => table_out <= 2983;
			WHEN "000110101101" => table_out <= 2984;
			WHEN "000110101110" => table_out <= 2985;
			WHEN "000110101111" => table_out <= 2986;
			WHEN "000110110000" => table_out <= 2987;
			WHEN "000110110001" => table_out <= 2989;
			WHEN "000110110010" => table_out <= 2990;
			WHEN "000110110011" => table_out <= 2991;
			WHEN "000110110100" => table_out <= 2992;
			WHEN "000110110101" => table_out <= 2993;
			WHEN "000110110110" => table_out <= 2994;
			WHEN "000110110111" => table_out <= 2995;
			WHEN "000110111000" => table_out <= 2996;
			WHEN "000110111001" => table_out <= 2998;
			WHEN "000110111010" => table_out <= 2999;
			WHEN "000110111011" => table_out <= 3000;
			WHEN "000110111100" => table_out <= 3001;
			WHEN "000110111101" => table_out <= 3002;
			WHEN "000110111110" => table_out <= 3003;
			WHEN "000110111111" => table_out <= 3004;
			WHEN "000111000000" => table_out <= 3005;
			WHEN "000111000001" => table_out <= 3006;
			WHEN "000111000010" => table_out <= 3008;
			WHEN "000111000011" => table_out <= 3009;
			WHEN "000111000100" => table_out <= 3010;
			WHEN "000111000101" => table_out <= 3011;
			WHEN "000111000110" => table_out <= 3012;
			WHEN "000111000111" => table_out <= 3013;
			WHEN "000111001000" => table_out <= 3014;
			WHEN "000111001001" => table_out <= 3015;
			WHEN "000111001010" => table_out <= 3016;
			WHEN "000111001011" => table_out <= 3017;
			WHEN "000111001100" => table_out <= 3018;
			WHEN "000111001101" => table_out <= 3019;
			WHEN "000111001110" => table_out <= 3021;
			WHEN "000111001111" => table_out <= 3022;
			WHEN "000111010000" => table_out <= 3023;
			WHEN "000111010001" => table_out <= 3024;
			WHEN "000111010010" => table_out <= 3025;
			WHEN "000111010011" => table_out <= 3026;
			WHEN "000111010100" => table_out <= 3027;
			WHEN "000111010101" => table_out <= 3028;
			WHEN "000111010110" => table_out <= 3029;
			WHEN "000111010111" => table_out <= 3030;
			WHEN "000111011000" => table_out <= 3031;
			WHEN "000111011001" => table_out <= 3032;
			WHEN "000111011010" => table_out <= 3033;
			WHEN "000111011011" => table_out <= 3034;
			WHEN "000111011100" => table_out <= 3035;
			WHEN "000111011101" => table_out <= 3036;
			WHEN "000111011110" => table_out <= 3037;
			WHEN "000111011111" => table_out <= 3038;
			WHEN "000111100000" => table_out <= 3039;
			WHEN "000111100001" => table_out <= 3040;
			WHEN "000111100010" => table_out <= 3041;
			WHEN "000111100011" => table_out <= 3042;
			WHEN "000111100100" => table_out <= 3043;
			WHEN "000111100101" => table_out <= 3044;
			WHEN "000111100110" => table_out <= 3045;
			WHEN "000111100111" => table_out <= 3046;
			WHEN "000111101000" => table_out <= 3047;
			WHEN "000111101001" => table_out <= 3048;
			WHEN "000111101010" => table_out <= 3049;
			WHEN "000111101011" => table_out <= 3050;
			WHEN "000111101100" => table_out <= 3051;
			WHEN "000111101101" => table_out <= 3052;
			WHEN "000111101110" => table_out <= 3053;
			WHEN "000111101111" => table_out <= 3054;
			WHEN "000111110000" => table_out <= 3055;
			WHEN "000111110001" => table_out <= 3056;
			WHEN "000111110010" => table_out <= 3057;
			WHEN "000111110011" => table_out <= 3058;
			WHEN "000111110100" => table_out <= 3059;
			WHEN "000111110101" => table_out <= 3060;
			WHEN "000111110110" => table_out <= 3061;
			WHEN "000111110111" => table_out <= 3062;
			WHEN "000111111000" => table_out <= 3063;
			WHEN "000111111001" => table_out <= 3064;
			WHEN "000111111010" => table_out <= 3065;
			WHEN "000111111011" => table_out <= 3066;
			WHEN "000111111100" => table_out <= 3067;
			WHEN "000111111101" => table_out <= 3068;
			WHEN "000111111110" => table_out <= 3069;
			WHEN "000111111111" => table_out <= 3070;
			WHEN "001000000000" => table_out <= 3071;
			WHEN "001000000001" => table_out <= 3072;
			WHEN "001000000010" => table_out <= 3073;
			WHEN "001000000011" => table_out <= 3074;
			WHEN "001000000100" => table_out <= 3075;
			WHEN "001000000101" => table_out <= 3076;
			WHEN "001000000110" => table_out <= 3077;
			WHEN "001000000111" => table_out <= 3078;
			WHEN "001000001000" => table_out <= 3079;
			WHEN "001000001001" => table_out <= 3080;
			WHEN "001000001010" => table_out <= 3081;
			WHEN "001000001011" => table_out <= 3082;
			WHEN "001000001100" => table_out <= 3082;
			WHEN "001000001101" => table_out <= 3083;
			WHEN "001000001110" => table_out <= 3084;
			WHEN "001000001111" => table_out <= 3085;
			WHEN "001000010000" => table_out <= 3086;
			WHEN "001000010001" => table_out <= 3087;
			WHEN "001000010010" => table_out <= 3088;
			WHEN "001000010011" => table_out <= 3089;
			WHEN "001000010100" => table_out <= 3090;
			WHEN "001000010101" => table_out <= 3091;
			WHEN "001000010110" => table_out <= 3092;
			WHEN "001000010111" => table_out <= 3093;
			WHEN "001000011000" => table_out <= 3094;
			WHEN "001000011001" => table_out <= 3095;
			WHEN "001000011010" => table_out <= 3095;
			WHEN "001000011011" => table_out <= 3096;
			WHEN "001000011100" => table_out <= 3097;
			WHEN "001000011101" => table_out <= 3098;
			WHEN "001000011110" => table_out <= 3099;
			WHEN "001000011111" => table_out <= 3100;
			WHEN "001000100000" => table_out <= 3101;
			WHEN "001000100001" => table_out <= 3102;
			WHEN "001000100010" => table_out <= 3103;
			WHEN "001000100011" => table_out <= 3104;
			WHEN "001000100100" => table_out <= 3105;
			WHEN "001000100101" => table_out <= 3105;
			WHEN "001000100110" => table_out <= 3106;
			WHEN "001000100111" => table_out <= 3107;
			WHEN "001000101000" => table_out <= 3108;
			WHEN "001000101001" => table_out <= 3109;
			WHEN "001000101010" => table_out <= 3110;
			WHEN "001000101011" => table_out <= 3111;
			WHEN "001000101100" => table_out <= 3112;
			WHEN "001000101101" => table_out <= 3113;
			WHEN "001000101110" => table_out <= 3113;
			WHEN "001000101111" => table_out <= 3114;
			WHEN "001000110000" => table_out <= 3115;
			WHEN "001000110001" => table_out <= 3116;
			WHEN "001000110010" => table_out <= 3117;
			WHEN "001000110011" => table_out <= 3118;
			WHEN "001000110100" => table_out <= 3119;
			WHEN "001000110101" => table_out <= 3120;
			WHEN "001000110110" => table_out <= 3120;
			WHEN "001000110111" => table_out <= 3121;
			WHEN "001000111000" => table_out <= 3122;
			WHEN "001000111001" => table_out <= 3123;
			WHEN "001000111010" => table_out <= 3124;
			WHEN "001000111011" => table_out <= 3125;
			WHEN "001000111100" => table_out <= 3126;
			WHEN "001000111101" => table_out <= 3126;
			WHEN "001000111110" => table_out <= 3127;
			WHEN "001000111111" => table_out <= 3128;
			WHEN "001001000000" => table_out <= 3129;
			WHEN "001001000001" => table_out <= 3130;
			WHEN "001001000010" => table_out <= 3131;
			WHEN "001001000011" => table_out <= 3132;
			WHEN "001001000100" => table_out <= 3132;
			WHEN "001001000101" => table_out <= 3133;
			WHEN "001001000110" => table_out <= 3134;
			WHEN "001001000111" => table_out <= 3135;
			WHEN "001001001000" => table_out <= 3136;
			WHEN "001001001001" => table_out <= 3137;
			WHEN "001001001010" => table_out <= 3138;
			WHEN "001001001011" => table_out <= 3138;
			WHEN "001001001100" => table_out <= 3139;
			WHEN "001001001101" => table_out <= 3140;
			WHEN "001001001110" => table_out <= 3141;
			WHEN "001001001111" => table_out <= 3142;
			WHEN "001001010000" => table_out <= 3143;
			WHEN "001001010001" => table_out <= 3143;
			WHEN "001001010010" => table_out <= 3144;
			WHEN "001001010011" => table_out <= 3145;
			WHEN "001001010100" => table_out <= 3146;
			WHEN "001001010101" => table_out <= 3147;
			WHEN "001001010110" => table_out <= 3148;
			WHEN "001001010111" => table_out <= 3148;
			WHEN "001001011000" => table_out <= 3149;
			WHEN "001001011001" => table_out <= 3150;
			WHEN "001001011010" => table_out <= 3151;
			WHEN "001001011011" => table_out <= 3152;
			WHEN "001001011100" => table_out <= 3152;
			WHEN "001001011101" => table_out <= 3153;
			WHEN "001001011110" => table_out <= 3154;
			WHEN "001001011111" => table_out <= 3155;
			WHEN "001001100000" => table_out <= 3156;
			WHEN "001001100001" => table_out <= 3156;
			WHEN "001001100010" => table_out <= 3157;
			WHEN "001001100011" => table_out <= 3158;
			WHEN "001001100100" => table_out <= 3159;
			WHEN "001001100101" => table_out <= 3160;
			WHEN "001001100110" => table_out <= 3161;
			WHEN "001001100111" => table_out <= 3161;
			WHEN "001001101000" => table_out <= 3162;
			WHEN "001001101001" => table_out <= 3163;
			WHEN "001001101010" => table_out <= 3164;
			WHEN "001001101011" => table_out <= 3165;
			WHEN "001001101100" => table_out <= 3165;
			WHEN "001001101101" => table_out <= 3166;
			WHEN "001001101110" => table_out <= 3167;
			WHEN "001001101111" => table_out <= 3168;
			WHEN "001001110000" => table_out <= 3168;
			WHEN "001001110001" => table_out <= 3169;
			WHEN "001001110010" => table_out <= 3170;
			WHEN "001001110011" => table_out <= 3171;
			WHEN "001001110100" => table_out <= 3172;
			WHEN "001001110101" => table_out <= 3172;
			WHEN "001001110110" => table_out <= 3173;
			WHEN "001001110111" => table_out <= 3174;
			WHEN "001001111000" => table_out <= 3175;
			WHEN "001001111001" => table_out <= 3176;
			WHEN "001001111010" => table_out <= 3176;
			WHEN "001001111011" => table_out <= 3177;
			WHEN "001001111100" => table_out <= 3178;
			WHEN "001001111101" => table_out <= 3179;
			WHEN "001001111110" => table_out <= 3179;
			WHEN "001001111111" => table_out <= 3180;
			WHEN "001010000000" => table_out <= 3181;
			WHEN "001010000001" => table_out <= 3182;
			WHEN "001010000010" => table_out <= 3182;
			WHEN "001010000011" => table_out <= 3183;
			WHEN "001010000100" => table_out <= 3184;
			WHEN "001010000101" => table_out <= 3185;
			WHEN "001010000110" => table_out <= 3186;
			WHEN "001010000111" => table_out <= 3186;
			WHEN "001010001000" => table_out <= 3187;
			WHEN "001010001001" => table_out <= 3188;
			WHEN "001010001010" => table_out <= 3189;
			WHEN "001010001011" => table_out <= 3189;
			WHEN "001010001100" => table_out <= 3190;
			WHEN "001010001101" => table_out <= 3191;
			WHEN "001010001110" => table_out <= 3192;
			WHEN "001010001111" => table_out <= 3192;
			WHEN "001010010000" => table_out <= 3193;
			WHEN "001010010001" => table_out <= 3194;
			WHEN "001010010010" => table_out <= 3195;
			WHEN "001010010011" => table_out <= 3195;
			WHEN "001010010100" => table_out <= 3196;
			WHEN "001010010101" => table_out <= 3197;
			WHEN "001010010110" => table_out <= 3198;
			WHEN "001010010111" => table_out <= 3198;
			WHEN "001010011000" => table_out <= 3199;
			WHEN "001010011001" => table_out <= 3200;
			WHEN "001010011010" => table_out <= 3201;
			WHEN "001010011011" => table_out <= 3201;
			WHEN "001010011100" => table_out <= 3202;
			WHEN "001010011101" => table_out <= 3203;
			WHEN "001010011110" => table_out <= 3203;
			WHEN "001010011111" => table_out <= 3204;
			WHEN "001010100000" => table_out <= 3205;
			WHEN "001010100001" => table_out <= 3206;
			WHEN "001010100010" => table_out <= 3206;
			WHEN "001010100011" => table_out <= 3207;
			WHEN "001010100100" => table_out <= 3208;
			WHEN "001010100101" => table_out <= 3209;
			WHEN "001010100110" => table_out <= 3209;
			WHEN "001010100111" => table_out <= 3210;
			WHEN "001010101000" => table_out <= 3211;
			WHEN "001010101001" => table_out <= 3211;
			WHEN "001010101010" => table_out <= 3212;
			WHEN "001010101011" => table_out <= 3213;
			WHEN "001010101100" => table_out <= 3214;
			WHEN "001010101101" => table_out <= 3214;
			WHEN "001010101110" => table_out <= 3215;
			WHEN "001010101111" => table_out <= 3216;
			WHEN "001010110000" => table_out <= 3217;
			WHEN "001010110001" => table_out <= 3217;
			WHEN "001010110010" => table_out <= 3218;
			WHEN "001010110011" => table_out <= 3219;
			WHEN "001010110100" => table_out <= 3219;
			WHEN "001010110101" => table_out <= 3220;
			WHEN "001010110110" => table_out <= 3221;
			WHEN "001010110111" => table_out <= 3222;
			WHEN "001010111000" => table_out <= 3222;
			WHEN "001010111001" => table_out <= 3223;
			WHEN "001010111010" => table_out <= 3224;
			WHEN "001010111011" => table_out <= 3224;
			WHEN "001010111100" => table_out <= 3225;
			WHEN "001010111101" => table_out <= 3226;
			WHEN "001010111110" => table_out <= 3226;
			WHEN "001010111111" => table_out <= 3227;
			WHEN "001011000000" => table_out <= 3228;
			WHEN "001011000001" => table_out <= 3229;
			WHEN "001011000010" => table_out <= 3229;
			WHEN "001011000011" => table_out <= 3230;
			WHEN "001011000100" => table_out <= 3231;
			WHEN "001011000101" => table_out <= 3231;
			WHEN "001011000110" => table_out <= 3232;
			WHEN "001011000111" => table_out <= 3233;
			WHEN "001011001000" => table_out <= 3233;
			WHEN "001011001001" => table_out <= 3234;
			WHEN "001011001010" => table_out <= 3235;
			WHEN "001011001011" => table_out <= 3235;
			WHEN "001011001100" => table_out <= 3236;
			WHEN "001011001101" => table_out <= 3237;
			WHEN "001011001110" => table_out <= 3238;
			WHEN "001011001111" => table_out <= 3238;
			WHEN "001011010000" => table_out <= 3239;
			WHEN "001011010001" => table_out <= 3240;
			WHEN "001011010010" => table_out <= 3240;
			WHEN "001011010011" => table_out <= 3241;
			WHEN "001011010100" => table_out <= 3242;
			WHEN "001011010101" => table_out <= 3242;
			WHEN "001011010110" => table_out <= 3243;
			WHEN "001011010111" => table_out <= 3244;
			WHEN "001011011000" => table_out <= 3244;
			WHEN "001011011001" => table_out <= 3245;
			WHEN "001011011010" => table_out <= 3246;
			WHEN "001011011011" => table_out <= 3246;
			WHEN "001011011100" => table_out <= 3247;
			WHEN "001011011101" => table_out <= 3248;
			WHEN "001011011110" => table_out <= 3248;
			WHEN "001011011111" => table_out <= 3249;
			WHEN "001011100000" => table_out <= 3250;
			WHEN "001011100001" => table_out <= 3250;
			WHEN "001011100010" => table_out <= 3251;
			WHEN "001011100011" => table_out <= 3252;
			WHEN "001011100100" => table_out <= 3252;
			WHEN "001011100101" => table_out <= 3253;
			WHEN "001011100110" => table_out <= 3254;
			WHEN "001011100111" => table_out <= 3254;
			WHEN "001011101000" => table_out <= 3255;
			WHEN "001011101001" => table_out <= 3256;
			WHEN "001011101010" => table_out <= 3256;
			WHEN "001011101011" => table_out <= 3257;
			WHEN "001011101100" => table_out <= 3258;
			WHEN "001011101101" => table_out <= 3258;
			WHEN "001011101110" => table_out <= 3259;
			WHEN "001011101111" => table_out <= 3260;
			WHEN "001011110000" => table_out <= 3260;
			WHEN "001011110001" => table_out <= 3261;
			WHEN "001011110010" => table_out <= 3262;
			WHEN "001011110011" => table_out <= 3262;
			WHEN "001011110100" => table_out <= 3263;
			WHEN "001011110101" => table_out <= 3264;
			WHEN "001011110110" => table_out <= 3264;
			WHEN "001011110111" => table_out <= 3265;
			WHEN "001011111000" => table_out <= 3266;
			WHEN "001011111001" => table_out <= 3266;
			WHEN "001011111010" => table_out <= 3267;
			WHEN "001011111011" => table_out <= 3267;
			WHEN "001011111100" => table_out <= 3268;
			WHEN "001011111101" => table_out <= 3269;
			WHEN "001011111110" => table_out <= 3269;
			WHEN "001011111111" => table_out <= 3270;
			WHEN "001100000000" => table_out <= 3271;
			WHEN "001100000001" => table_out <= 3271;
			WHEN "001100000010" => table_out <= 3272;
			WHEN "001100000011" => table_out <= 3273;
			WHEN "001100000100" => table_out <= 3273;
			WHEN "001100000101" => table_out <= 3274;
			WHEN "001100000110" => table_out <= 3274;
			WHEN "001100000111" => table_out <= 3275;
			WHEN "001100001000" => table_out <= 3276;
			WHEN "001100001001" => table_out <= 3276;
			WHEN "001100001010" => table_out <= 3277;
			WHEN "001100001011" => table_out <= 3278;
			WHEN "001100001100" => table_out <= 3278;
			WHEN "001100001101" => table_out <= 3279;
			WHEN "001100001110" => table_out <= 3280;
			WHEN "001100001111" => table_out <= 3280;
			WHEN "001100010000" => table_out <= 3281;
			WHEN "001100010001" => table_out <= 3281;
			WHEN "001100010010" => table_out <= 3282;
			WHEN "001100010011" => table_out <= 3283;
			WHEN "001100010100" => table_out <= 3283;
			WHEN "001100010101" => table_out <= 3284;
			WHEN "001100010110" => table_out <= 3285;
			WHEN "001100010111" => table_out <= 3285;
			WHEN "001100011000" => table_out <= 3286;
			WHEN "001100011001" => table_out <= 3286;
			WHEN "001100011010" => table_out <= 3287;
			WHEN "001100011011" => table_out <= 3288;
			WHEN "001100011100" => table_out <= 3288;
			WHEN "001100011101" => table_out <= 3289;
			WHEN "001100011110" => table_out <= 3290;
			WHEN "001100011111" => table_out <= 3290;
			WHEN "001100100000" => table_out <= 3291;
			WHEN "001100100001" => table_out <= 3291;
			WHEN "001100100010" => table_out <= 3292;
			WHEN "001100100011" => table_out <= 3293;
			WHEN "001100100100" => table_out <= 3293;
			WHEN "001100100101" => table_out <= 3294;
			WHEN "001100100110" => table_out <= 3294;
			WHEN "001100100111" => table_out <= 3295;
			WHEN "001100101000" => table_out <= 3296;
			WHEN "001100101001" => table_out <= 3296;
			WHEN "001100101010" => table_out <= 3297;
			WHEN "001100101011" => table_out <= 3297;
			WHEN "001100101100" => table_out <= 3298;
			WHEN "001100101101" => table_out <= 3299;
			WHEN "001100101110" => table_out <= 3299;
			WHEN "001100101111" => table_out <= 3300;
			WHEN "001100110000" => table_out <= 3301;
			WHEN "001100110001" => table_out <= 3301;
			WHEN "001100110010" => table_out <= 3302;
			WHEN "001100110011" => table_out <= 3302;
			WHEN "001100110100" => table_out <= 3303;
			WHEN "001100110101" => table_out <= 3304;
			WHEN "001100110110" => table_out <= 3304;
			WHEN "001100110111" => table_out <= 3305;
			WHEN "001100111000" => table_out <= 3305;
			WHEN "001100111001" => table_out <= 3306;
			WHEN "001100111010" => table_out <= 3307;
			WHEN "001100111011" => table_out <= 3307;
			WHEN "001100111100" => table_out <= 3308;
			WHEN "001100111101" => table_out <= 3308;
			WHEN "001100111110" => table_out <= 3309;
			WHEN "001100111111" => table_out <= 3309;
			WHEN "001101000000" => table_out <= 3310;
			WHEN "001101000001" => table_out <= 3311;
			WHEN "001101000010" => table_out <= 3311;
			WHEN "001101000011" => table_out <= 3312;
			WHEN "001101000100" => table_out <= 3312;
			WHEN "001101000101" => table_out <= 3313;
			WHEN "001101000110" => table_out <= 3314;
			WHEN "001101000111" => table_out <= 3314;
			WHEN "001101001000" => table_out <= 3315;
			WHEN "001101001001" => table_out <= 3315;
			WHEN "001101001010" => table_out <= 3316;
			WHEN "001101001011" => table_out <= 3317;
			WHEN "001101001100" => table_out <= 3317;
			WHEN "001101001101" => table_out <= 3318;
			WHEN "001101001110" => table_out <= 3318;
			WHEN "001101001111" => table_out <= 3319;
			WHEN "001101010000" => table_out <= 3319;
			WHEN "001101010001" => table_out <= 3320;
			WHEN "001101010010" => table_out <= 3321;
			WHEN "001101010011" => table_out <= 3321;
			WHEN "001101010100" => table_out <= 3322;
			WHEN "001101010101" => table_out <= 3322;
			WHEN "001101010110" => table_out <= 3323;
			WHEN "001101010111" => table_out <= 3323;
			WHEN "001101011000" => table_out <= 3324;
			WHEN "001101011001" => table_out <= 3325;
			WHEN "001101011010" => table_out <= 3325;
			WHEN "001101011011" => table_out <= 3326;
			WHEN "001101011100" => table_out <= 3326;
			WHEN "001101011101" => table_out <= 3327;
			WHEN "001101011110" => table_out <= 3327;
			WHEN "001101011111" => table_out <= 3328;
			WHEN "001101100000" => table_out <= 3329;
			WHEN "001101100001" => table_out <= 3329;
			WHEN "001101100010" => table_out <= 3330;
			WHEN "001101100011" => table_out <= 3330;
			WHEN "001101100100" => table_out <= 3331;
			WHEN "001101100101" => table_out <= 3331;
			WHEN "001101100110" => table_out <= 3332;
			WHEN "001101100111" => table_out <= 3333;
			WHEN "001101101000" => table_out <= 3333;
			WHEN "001101101001" => table_out <= 3334;
			WHEN "001101101010" => table_out <= 3334;
			WHEN "001101101011" => table_out <= 3335;
			WHEN "001101101100" => table_out <= 3335;
			WHEN "001101101101" => table_out <= 3336;
			WHEN "001101101110" => table_out <= 3337;
			WHEN "001101101111" => table_out <= 3337;
			WHEN "001101110000" => table_out <= 3338;
			WHEN "001101110001" => table_out <= 3338;
			WHEN "001101110010" => table_out <= 3339;
			WHEN "001101110011" => table_out <= 3339;
			WHEN "001101110100" => table_out <= 3340;
			WHEN "001101110101" => table_out <= 3340;
			WHEN "001101110110" => table_out <= 3341;
			WHEN "001101110111" => table_out <= 3342;
			WHEN "001101111000" => table_out <= 3342;
			WHEN "001101111001" => table_out <= 3343;
			WHEN "001101111010" => table_out <= 3343;
			WHEN "001101111011" => table_out <= 3344;
			WHEN "001101111100" => table_out <= 3344;
			WHEN "001101111101" => table_out <= 3345;
			WHEN "001101111110" => table_out <= 3345;
			WHEN "001101111111" => table_out <= 3346;
			WHEN "001110000000" => table_out <= 3347;
			WHEN "001110000001" => table_out <= 3347;
			WHEN "001110000010" => table_out <= 3348;
			WHEN "001110000011" => table_out <= 3348;
			WHEN "001110000100" => table_out <= 3349;
			WHEN "001110000101" => table_out <= 3349;
			WHEN "001110000110" => table_out <= 3350;
			WHEN "001110000111" => table_out <= 3350;
			WHEN "001110001000" => table_out <= 3351;
			WHEN "001110001001" => table_out <= 3351;
			WHEN "001110001010" => table_out <= 3352;
			WHEN "001110001011" => table_out <= 3353;
			WHEN "001110001100" => table_out <= 3353;
			WHEN "001110001101" => table_out <= 3354;
			WHEN "001110001110" => table_out <= 3354;
			WHEN "001110001111" => table_out <= 3355;
			WHEN "001110010000" => table_out <= 3355;
			WHEN "001110010001" => table_out <= 3356;
			WHEN "001110010010" => table_out <= 3356;
			WHEN "001110010011" => table_out <= 3357;
			WHEN "001110010100" => table_out <= 3357;
			WHEN "001110010101" => table_out <= 3358;
			WHEN "001110010110" => table_out <= 3358;
			WHEN "001110010111" => table_out <= 3359;
			WHEN "001110011000" => table_out <= 3360;
			WHEN "001110011001" => table_out <= 3360;
			WHEN "001110011010" => table_out <= 3361;
			WHEN "001110011011" => table_out <= 3361;
			WHEN "001110011100" => table_out <= 3362;
			WHEN "001110011101" => table_out <= 3362;
			WHEN "001110011110" => table_out <= 3363;
			WHEN "001110011111" => table_out <= 3363;
			WHEN "001110100000" => table_out <= 3364;
			WHEN "001110100001" => table_out <= 3364;
			WHEN "001110100010" => table_out <= 3365;
			WHEN "001110100011" => table_out <= 3365;
			WHEN "001110100100" => table_out <= 3366;
			WHEN "001110100101" => table_out <= 3366;
			WHEN "001110100110" => table_out <= 3367;
			WHEN "001110100111" => table_out <= 3368;
			WHEN "001110101000" => table_out <= 3368;
			WHEN "001110101001" => table_out <= 3369;
			WHEN "001110101010" => table_out <= 3369;
			WHEN "001110101011" => table_out <= 3370;
			WHEN "001110101100" => table_out <= 3370;
			WHEN "001110101101" => table_out <= 3371;
			WHEN "001110101110" => table_out <= 3371;
			WHEN "001110101111" => table_out <= 3372;
			WHEN "001110110000" => table_out <= 3372;
			WHEN "001110110001" => table_out <= 3373;
			WHEN "001110110010" => table_out <= 3373;
			WHEN "001110110011" => table_out <= 3374;
			WHEN "001110110100" => table_out <= 3374;
			WHEN "001110110101" => table_out <= 3375;
			WHEN "001110110110" => table_out <= 3375;
			WHEN "001110110111" => table_out <= 3376;
			WHEN "001110111000" => table_out <= 3376;
			WHEN "001110111001" => table_out <= 3377;
			WHEN "001110111010" => table_out <= 3377;
			WHEN "001110111011" => table_out <= 3378;
			WHEN "001110111100" => table_out <= 3378;
			WHEN "001110111101" => table_out <= 3379;
			WHEN "001110111110" => table_out <= 3379;
			WHEN "001110111111" => table_out <= 3380;
			WHEN "001111000000" => table_out <= 3381;
			WHEN "001111000001" => table_out <= 3381;
			WHEN "001111000010" => table_out <= 3382;
			WHEN "001111000011" => table_out <= 3382;
			WHEN "001111000100" => table_out <= 3383;
			WHEN "001111000101" => table_out <= 3383;
			WHEN "001111000110" => table_out <= 3384;
			WHEN "001111000111" => table_out <= 3384;
			WHEN "001111001000" => table_out <= 3385;
			WHEN "001111001001" => table_out <= 3385;
			WHEN "001111001010" => table_out <= 3386;
			WHEN "001111001011" => table_out <= 3386;
			WHEN "001111001100" => table_out <= 3387;
			WHEN "001111001101" => table_out <= 3387;
			WHEN "001111001110" => table_out <= 3388;
			WHEN "001111001111" => table_out <= 3388;
			WHEN "001111010000" => table_out <= 3389;
			WHEN "001111010001" => table_out <= 3389;
			WHEN "001111010010" => table_out <= 3390;
			WHEN "001111010011" => table_out <= 3390;
			WHEN "001111010100" => table_out <= 3391;
			WHEN "001111010101" => table_out <= 3391;
			WHEN "001111010110" => table_out <= 3392;
			WHEN "001111010111" => table_out <= 3392;
			WHEN "001111011000" => table_out <= 3393;
			WHEN "001111011001" => table_out <= 3393;
			WHEN "001111011010" => table_out <= 3394;
			WHEN "001111011011" => table_out <= 3394;
			WHEN "001111011100" => table_out <= 3395;
			WHEN "001111011101" => table_out <= 3395;
			WHEN "001111011110" => table_out <= 3396;
			WHEN "001111011111" => table_out <= 3396;
			WHEN "001111100000" => table_out <= 3397;
			WHEN "001111100001" => table_out <= 3397;
			WHEN "001111100010" => table_out <= 3398;
			WHEN "001111100011" => table_out <= 3398;
			WHEN "001111100100" => table_out <= 3399;
			WHEN "001111100101" => table_out <= 3399;
			WHEN "001111100110" => table_out <= 3400;
			WHEN "001111100111" => table_out <= 3400;
			WHEN "001111101000" => table_out <= 3401;
			WHEN "001111101001" => table_out <= 3401;
			WHEN "001111101010" => table_out <= 3402;
			WHEN "001111101011" => table_out <= 3402;
			WHEN "001111101100" => table_out <= 3403;
			WHEN "001111101101" => table_out <= 3403;
			WHEN "001111101110" => table_out <= 3404;
			WHEN "001111101111" => table_out <= 3404;
			WHEN "001111110000" => table_out <= 3405;
			WHEN "001111110001" => table_out <= 3405;
			WHEN "001111110010" => table_out <= 3405;
			WHEN "001111110011" => table_out <= 3406;
			WHEN "001111110100" => table_out <= 3406;
			WHEN "001111110101" => table_out <= 3407;
			WHEN "001111110110" => table_out <= 3407;
			WHEN "001111110111" => table_out <= 3408;
			WHEN "001111111000" => table_out <= 3408;
			WHEN "001111111001" => table_out <= 3409;
			WHEN "001111111010" => table_out <= 3409;
			WHEN "001111111011" => table_out <= 3410;
			WHEN "001111111100" => table_out <= 3410;
			WHEN "001111111101" => table_out <= 3411;
			WHEN "001111111110" => table_out <= 3411;
			WHEN "001111111111" => table_out <= 3412;
			WHEN "010000000000" => table_out <= 3412;
			WHEN "010000000001" => table_out <= 3413;
			WHEN "010000000010" => table_out <= 3413;
			WHEN "010000000011" => table_out <= 3414;
			WHEN "010000000100" => table_out <= 3414;
			WHEN "010000000101" => table_out <= 3415;
			WHEN "010000000110" => table_out <= 3415;
			WHEN "010000000111" => table_out <= 3416;
			WHEN "010000001000" => table_out <= 3416;
			WHEN "010000001001" => table_out <= 3417;
			WHEN "010000001010" => table_out <= 3417;
			WHEN "010000001011" => table_out <= 3418;
			WHEN "010000001100" => table_out <= 3418;
			WHEN "010000001101" => table_out <= 3418;
			WHEN "010000001110" => table_out <= 3419;
			WHEN "010000001111" => table_out <= 3419;
			WHEN "010000010000" => table_out <= 3420;
			WHEN "010000010001" => table_out <= 3420;
			WHEN "010000010010" => table_out <= 3421;
			WHEN "010000010011" => table_out <= 3421;
			WHEN "010000010100" => table_out <= 3422;
			WHEN "010000010101" => table_out <= 3422;
			WHEN "010000010110" => table_out <= 3423;
			WHEN "010000010111" => table_out <= 3423;
			WHEN "010000011000" => table_out <= 3424;
			WHEN "010000011001" => table_out <= 3424;
			WHEN "010000011010" => table_out <= 3425;
			WHEN "010000011011" => table_out <= 3425;
			WHEN "010000011100" => table_out <= 3426;
			WHEN "010000011101" => table_out <= 3426;
			WHEN "010000011110" => table_out <= 3426;
			WHEN "010000011111" => table_out <= 3427;
			WHEN "010000100000" => table_out <= 3427;
			WHEN "010000100001" => table_out <= 3428;
			WHEN "010000100010" => table_out <= 3428;
			WHEN "010000100011" => table_out <= 3429;
			WHEN "010000100100" => table_out <= 3429;
			WHEN "010000100101" => table_out <= 3430;
			WHEN "010000100110" => table_out <= 3430;
			WHEN "010000100111" => table_out <= 3431;
			WHEN "010000101000" => table_out <= 3431;
			WHEN "010000101001" => table_out <= 3432;
			WHEN "010000101010" => table_out <= 3432;
			WHEN "010000101011" => table_out <= 3433;
			WHEN "010000101100" => table_out <= 3433;
			WHEN "010000101101" => table_out <= 3433;
			WHEN "010000101110" => table_out <= 3434;
			WHEN "010000101111" => table_out <= 3434;
			WHEN "010000110000" => table_out <= 3435;
			WHEN "010000110001" => table_out <= 3435;
			WHEN "010000110010" => table_out <= 3436;
			WHEN "010000110011" => table_out <= 3436;
			WHEN "010000110100" => table_out <= 3437;
			WHEN "010000110101" => table_out <= 3437;
			WHEN "010000110110" => table_out <= 3438;
			WHEN "010000110111" => table_out <= 3438;
			WHEN "010000111000" => table_out <= 3438;
			WHEN "010000111001" => table_out <= 3439;
			WHEN "010000111010" => table_out <= 3439;
			WHEN "010000111011" => table_out <= 3440;
			WHEN "010000111100" => table_out <= 3440;
			WHEN "010000111101" => table_out <= 3441;
			WHEN "010000111110" => table_out <= 3441;
			WHEN "010000111111" => table_out <= 3442;
			WHEN "010001000000" => table_out <= 3442;
			WHEN "010001000001" => table_out <= 3443;
			WHEN "010001000010" => table_out <= 3443;
			WHEN "010001000011" => table_out <= 3443;
			WHEN "010001000100" => table_out <= 3444;
			WHEN "010001000101" => table_out <= 3444;
			WHEN "010001000110" => table_out <= 3445;
			WHEN "010001000111" => table_out <= 3445;
			WHEN "010001001000" => table_out <= 3446;
			WHEN "010001001001" => table_out <= 3446;
			WHEN "010001001010" => table_out <= 3447;
			WHEN "010001001011" => table_out <= 3447;
			WHEN "010001001100" => table_out <= 3448;
			WHEN "010001001101" => table_out <= 3448;
			WHEN "010001001110" => table_out <= 3448;
			WHEN "010001001111" => table_out <= 3449;
			WHEN "010001010000" => table_out <= 3449;
			WHEN "010001010001" => table_out <= 3450;
			WHEN "010001010010" => table_out <= 3450;
			WHEN "010001010011" => table_out <= 3451;
			WHEN "010001010100" => table_out <= 3451;
			WHEN "010001010101" => table_out <= 3452;
			WHEN "010001010110" => table_out <= 3452;
			WHEN "010001010111" => table_out <= 3452;
			WHEN "010001011000" => table_out <= 3453;
			WHEN "010001011001" => table_out <= 3453;
			WHEN "010001011010" => table_out <= 3454;
			WHEN "010001011011" => table_out <= 3454;
			WHEN "010001011100" => table_out <= 3455;
			WHEN "010001011101" => table_out <= 3455;
			WHEN "010001011110" => table_out <= 3455;
			WHEN "010001011111" => table_out <= 3456;
			WHEN "010001100000" => table_out <= 3456;
			WHEN "010001100001" => table_out <= 3457;
			WHEN "010001100010" => table_out <= 3457;
			WHEN "010001100011" => table_out <= 3458;
			WHEN "010001100100" => table_out <= 3458;
			WHEN "010001100101" => table_out <= 3459;
			WHEN "010001100110" => table_out <= 3459;
			WHEN "010001100111" => table_out <= 3459;
			WHEN "010001101000" => table_out <= 3460;
			WHEN "010001101001" => table_out <= 3460;
			WHEN "010001101010" => table_out <= 3461;
			WHEN "010001101011" => table_out <= 3461;
			WHEN "010001101100" => table_out <= 3462;
			WHEN "010001101101" => table_out <= 3462;
			WHEN "010001101110" => table_out <= 3462;
			WHEN "010001101111" => table_out <= 3463;
			WHEN "010001110000" => table_out <= 3463;
			WHEN "010001110001" => table_out <= 3464;
			WHEN "010001110010" => table_out <= 3464;
			WHEN "010001110011" => table_out <= 3465;
			WHEN "010001110100" => table_out <= 3465;
			WHEN "010001110101" => table_out <= 3466;
			WHEN "010001110110" => table_out <= 3466;
			WHEN "010001110111" => table_out <= 3466;
			WHEN "010001111000" => table_out <= 3467;
			WHEN "010001111001" => table_out <= 3467;
			WHEN "010001111010" => table_out <= 3468;
			WHEN "010001111011" => table_out <= 3468;
			WHEN "010001111100" => table_out <= 3469;
			WHEN "010001111101" => table_out <= 3469;
			WHEN "010001111110" => table_out <= 3469;
			WHEN "010001111111" => table_out <= 3470;
			WHEN "010010000000" => table_out <= 3470;
			WHEN "010010000001" => table_out <= 3471;
			WHEN "010010000010" => table_out <= 3471;
			WHEN "010010000011" => table_out <= 3472;
			WHEN "010010000100" => table_out <= 3472;
			WHEN "010010000101" => table_out <= 3472;
			WHEN "010010000110" => table_out <= 3473;
			WHEN "010010000111" => table_out <= 3473;
			WHEN "010010001000" => table_out <= 3474;
			WHEN "010010001001" => table_out <= 3474;
			WHEN "010010001010" => table_out <= 3474;
			WHEN "010010001011" => table_out <= 3475;
			WHEN "010010001100" => table_out <= 3475;
			WHEN "010010001101" => table_out <= 3476;
			WHEN "010010001110" => table_out <= 3476;
			WHEN "010010001111" => table_out <= 3477;
			WHEN "010010010000" => table_out <= 3477;
			WHEN "010010010001" => table_out <= 3477;
			WHEN "010010010010" => table_out <= 3478;
			WHEN "010010010011" => table_out <= 3478;
			WHEN "010010010100" => table_out <= 3479;
			WHEN "010010010101" => table_out <= 3479;
			WHEN "010010010110" => table_out <= 3480;
			WHEN "010010010111" => table_out <= 3480;
			WHEN "010010011000" => table_out <= 3480;
			WHEN "010010011001" => table_out <= 3481;
			WHEN "010010011010" => table_out <= 3481;
			WHEN "010010011011" => table_out <= 3482;
			WHEN "010010011100" => table_out <= 3482;
			WHEN "010010011101" => table_out <= 3482;
			WHEN "010010011110" => table_out <= 3483;
			WHEN "010010011111" => table_out <= 3483;
			WHEN "010010100000" => table_out <= 3484;
			WHEN "010010100001" => table_out <= 3484;
			WHEN "010010100010" => table_out <= 3485;
			WHEN "010010100011" => table_out <= 3485;
			WHEN "010010100100" => table_out <= 3485;
			WHEN "010010100101" => table_out <= 3486;
			WHEN "010010100110" => table_out <= 3486;
			WHEN "010010100111" => table_out <= 3487;
			WHEN "010010101000" => table_out <= 3487;
			WHEN "010010101001" => table_out <= 3487;
			WHEN "010010101010" => table_out <= 3488;
			WHEN "010010101011" => table_out <= 3488;
			WHEN "010010101100" => table_out <= 3489;
			WHEN "010010101101" => table_out <= 3489;
			WHEN "010010101110" => table_out <= 3490;
			WHEN "010010101111" => table_out <= 3490;
			WHEN "010010110000" => table_out <= 3490;
			WHEN "010010110001" => table_out <= 3491;
			WHEN "010010110010" => table_out <= 3491;
			WHEN "010010110011" => table_out <= 3492;
			WHEN "010010110100" => table_out <= 3492;
			WHEN "010010110101" => table_out <= 3492;
			WHEN "010010110110" => table_out <= 3493;
			WHEN "010010110111" => table_out <= 3493;
			WHEN "010010111000" => table_out <= 3494;
			WHEN "010010111001" => table_out <= 3494;
			WHEN "010010111010" => table_out <= 3494;
			WHEN "010010111011" => table_out <= 3495;
			WHEN "010010111100" => table_out <= 3495;
			WHEN "010010111101" => table_out <= 3496;
			WHEN "010010111110" => table_out <= 3496;
			WHEN "010010111111" => table_out <= 3496;
			WHEN "010011000000" => table_out <= 3497;
			WHEN "010011000001" => table_out <= 3497;
			WHEN "010011000010" => table_out <= 3498;
			WHEN "010011000011" => table_out <= 3498;
			WHEN "010011000100" => table_out <= 3498;
			WHEN "010011000101" => table_out <= 3499;
			WHEN "010011000110" => table_out <= 3499;
			WHEN "010011000111" => table_out <= 3500;
			WHEN "010011001000" => table_out <= 3500;
			WHEN "010011001001" => table_out <= 3500;
			WHEN "010011001010" => table_out <= 3501;
			WHEN "010011001011" => table_out <= 3501;
			WHEN "010011001100" => table_out <= 3502;
			WHEN "010011001101" => table_out <= 3502;
			WHEN "010011001110" => table_out <= 3502;
			WHEN "010011001111" => table_out <= 3503;
			WHEN "010011010000" => table_out <= 3503;
			WHEN "010011010001" => table_out <= 3504;
			WHEN "010011010010" => table_out <= 3504;
			WHEN "010011010011" => table_out <= 3504;
			WHEN "010011010100" => table_out <= 3505;
			WHEN "010011010101" => table_out <= 3505;
			WHEN "010011010110" => table_out <= 3506;
			WHEN "010011010111" => table_out <= 3506;
			WHEN "010011011000" => table_out <= 3506;
			WHEN "010011011001" => table_out <= 3507;
			WHEN "010011011010" => table_out <= 3507;
			WHEN "010011011011" => table_out <= 3508;
			WHEN "010011011100" => table_out <= 3508;
			WHEN "010011011101" => table_out <= 3508;
			WHEN "010011011110" => table_out <= 3509;
			WHEN "010011011111" => table_out <= 3509;
			WHEN "010011100000" => table_out <= 3510;
			WHEN "010011100001" => table_out <= 3510;
			WHEN "010011100010" => table_out <= 3510;
			WHEN "010011100011" => table_out <= 3511;
			WHEN "010011100100" => table_out <= 3511;
			WHEN "010011100101" => table_out <= 3512;
			WHEN "010011100110" => table_out <= 3512;
			WHEN "010011100111" => table_out <= 3512;
			WHEN "010011101000" => table_out <= 3513;
			WHEN "010011101001" => table_out <= 3513;
			WHEN "010011101010" => table_out <= 3514;
			WHEN "010011101011" => table_out <= 3514;
			WHEN "010011101100" => table_out <= 3514;
			WHEN "010011101101" => table_out <= 3515;
			WHEN "010011101110" => table_out <= 3515;
			WHEN "010011101111" => table_out <= 3516;
			WHEN "010011110000" => table_out <= 3516;
			WHEN "010011110001" => table_out <= 3516;
			WHEN "010011110010" => table_out <= 3517;
			WHEN "010011110011" => table_out <= 3517;
			WHEN "010011110100" => table_out <= 3517;
			WHEN "010011110101" => table_out <= 3518;
			WHEN "010011110110" => table_out <= 3518;
			WHEN "010011110111" => table_out <= 3519;
			WHEN "010011111000" => table_out <= 3519;
			WHEN "010011111001" => table_out <= 3519;
			WHEN "010011111010" => table_out <= 3520;
			WHEN "010011111011" => table_out <= 3520;
			WHEN "010011111100" => table_out <= 3521;
			WHEN "010011111101" => table_out <= 3521;
			WHEN "010011111110" => table_out <= 3521;
			WHEN "010011111111" => table_out <= 3522;
			WHEN "010100000000" => table_out <= 3522;
			WHEN "010100000001" => table_out <= 3522;
			WHEN "010100000010" => table_out <= 3523;
			WHEN "010100000011" => table_out <= 3523;
			WHEN "010100000100" => table_out <= 3524;
			WHEN "010100000101" => table_out <= 3524;
			WHEN "010100000110" => table_out <= 3524;
			WHEN "010100000111" => table_out <= 3525;
			WHEN "010100001000" => table_out <= 3525;
			WHEN "010100001001" => table_out <= 3526;
			WHEN "010100001010" => table_out <= 3526;
			WHEN "010100001011" => table_out <= 3526;
			WHEN "010100001100" => table_out <= 3527;
			WHEN "010100001101" => table_out <= 3527;
			WHEN "010100001110" => table_out <= 3527;
			WHEN "010100001111" => table_out <= 3528;
			WHEN "010100010000" => table_out <= 3528;
			WHEN "010100010001" => table_out <= 3529;
			WHEN "010100010010" => table_out <= 3529;
			WHEN "010100010011" => table_out <= 3529;
			WHEN "010100010100" => table_out <= 3530;
			WHEN "010100010101" => table_out <= 3530;
			WHEN "010100010110" => table_out <= 3530;
			WHEN "010100010111" => table_out <= 3531;
			WHEN "010100011000" => table_out <= 3531;
			WHEN "010100011001" => table_out <= 3532;
			WHEN "010100011010" => table_out <= 3532;
			WHEN "010100011011" => table_out <= 3532;
			WHEN "010100011100" => table_out <= 3533;
			WHEN "010100011101" => table_out <= 3533;
			WHEN "010100011110" => table_out <= 3534;
			WHEN "010100011111" => table_out <= 3534;
			WHEN "010100100000" => table_out <= 3534;
			WHEN "010100100001" => table_out <= 3535;
			WHEN "010100100010" => table_out <= 3535;
			WHEN "010100100011" => table_out <= 3535;
			WHEN "010100100100" => table_out <= 3536;
			WHEN "010100100101" => table_out <= 3536;
			WHEN "010100100110" => table_out <= 3537;
			WHEN "010100100111" => table_out <= 3537;
			WHEN "010100101000" => table_out <= 3537;
			WHEN "010100101001" => table_out <= 3538;
			WHEN "010100101010" => table_out <= 3538;
			WHEN "010100101011" => table_out <= 3538;
			WHEN "010100101100" => table_out <= 3539;
			WHEN "010100101101" => table_out <= 3539;
			WHEN "010100101110" => table_out <= 3539;
			WHEN "010100101111" => table_out <= 3540;
			WHEN "010100110000" => table_out <= 3540;
			WHEN "010100110001" => table_out <= 3541;
			WHEN "010100110010" => table_out <= 3541;
			WHEN "010100110011" => table_out <= 3541;
			WHEN "010100110100" => table_out <= 3542;
			WHEN "010100110101" => table_out <= 3542;
			WHEN "010100110110" => table_out <= 3542;
			WHEN "010100110111" => table_out <= 3543;
			WHEN "010100111000" => table_out <= 3543;
			WHEN "010100111001" => table_out <= 3544;
			WHEN "010100111010" => table_out <= 3544;
			WHEN "010100111011" => table_out <= 3544;
			WHEN "010100111100" => table_out <= 3545;
			WHEN "010100111101" => table_out <= 3545;
			WHEN "010100111110" => table_out <= 3545;
			WHEN "010100111111" => table_out <= 3546;
			WHEN "010101000000" => table_out <= 3546;
			WHEN "010101000001" => table_out <= 3546;
			WHEN "010101000010" => table_out <= 3547;
			WHEN "010101000011" => table_out <= 3547;
			WHEN "010101000100" => table_out <= 3548;
			WHEN "010101000101" => table_out <= 3548;
			WHEN "010101000110" => table_out <= 3548;
			WHEN "010101000111" => table_out <= 3549;
			WHEN "010101001000" => table_out <= 3549;
			WHEN "010101001001" => table_out <= 3549;
			WHEN "010101001010" => table_out <= 3550;
			WHEN "010101001011" => table_out <= 3550;
			WHEN "010101001100" => table_out <= 3550;
			WHEN "010101001101" => table_out <= 3551;
			WHEN "010101001110" => table_out <= 3551;
			WHEN "010101001111" => table_out <= 3552;
			WHEN "010101010000" => table_out <= 3552;
			WHEN "010101010001" => table_out <= 3552;
			WHEN "010101010010" => table_out <= 3553;
			WHEN "010101010011" => table_out <= 3553;
			WHEN "010101010100" => table_out <= 3553;
			WHEN "010101010101" => table_out <= 3554;
			WHEN "010101010110" => table_out <= 3554;
			WHEN "010101010111" => table_out <= 3554;
			WHEN "010101011000" => table_out <= 3555;
			WHEN "010101011001" => table_out <= 3555;
			WHEN "010101011010" => table_out <= 3556;
			WHEN "010101011011" => table_out <= 3556;
			WHEN "010101011100" => table_out <= 3556;
			WHEN "010101011101" => table_out <= 3557;
			WHEN "010101011110" => table_out <= 3557;
			WHEN "010101011111" => table_out <= 3557;
			WHEN "010101100000" => table_out <= 3558;
			WHEN "010101100001" => table_out <= 3558;
			WHEN "010101100010" => table_out <= 3558;
			WHEN "010101100011" => table_out <= 3559;
			WHEN "010101100100" => table_out <= 3559;
			WHEN "010101100101" => table_out <= 3559;
			WHEN "010101100110" => table_out <= 3560;
			WHEN "010101100111" => table_out <= 3560;
			WHEN "010101101000" => table_out <= 3561;
			WHEN "010101101001" => table_out <= 3561;
			WHEN "010101101010" => table_out <= 3561;
			WHEN "010101101011" => table_out <= 3562;
			WHEN "010101101100" => table_out <= 3562;
			WHEN "010101101101" => table_out <= 3562;
			WHEN "010101101110" => table_out <= 3563;
			WHEN "010101101111" => table_out <= 3563;
			WHEN "010101110000" => table_out <= 3563;
			WHEN "010101110001" => table_out <= 3564;
			WHEN "010101110010" => table_out <= 3564;
			WHEN "010101110011" => table_out <= 3564;
			WHEN "010101110100" => table_out <= 3565;
			WHEN "010101110101" => table_out <= 3565;
			WHEN "010101110110" => table_out <= 3566;
			WHEN "010101110111" => table_out <= 3566;
			WHEN "010101111000" => table_out <= 3566;
			WHEN "010101111001" => table_out <= 3567;
			WHEN "010101111010" => table_out <= 3567;
			WHEN "010101111011" => table_out <= 3567;
			WHEN "010101111100" => table_out <= 3568;
			WHEN "010101111101" => table_out <= 3568;
			WHEN "010101111110" => table_out <= 3568;
			WHEN "010101111111" => table_out <= 3569;
			WHEN "010110000000" => table_out <= 3569;
			WHEN "010110000001" => table_out <= 3569;
			WHEN "010110000010" => table_out <= 3570;
			WHEN "010110000011" => table_out <= 3570;
			WHEN "010110000100" => table_out <= 3570;
			WHEN "010110000101" => table_out <= 3571;
			WHEN "010110000110" => table_out <= 3571;
			WHEN "010110000111" => table_out <= 3571;
			WHEN "010110001000" => table_out <= 3572;
			WHEN "010110001001" => table_out <= 3572;
			WHEN "010110001010" => table_out <= 3572;
			WHEN "010110001011" => table_out <= 3573;
			WHEN "010110001100" => table_out <= 3573;
			WHEN "010110001101" => table_out <= 3574;
			WHEN "010110001110" => table_out <= 3574;
			WHEN "010110001111" => table_out <= 3574;
			WHEN "010110010000" => table_out <= 3575;
			WHEN "010110010001" => table_out <= 3575;
			WHEN "010110010010" => table_out <= 3575;
			WHEN "010110010011" => table_out <= 3576;
			WHEN "010110010100" => table_out <= 3576;
			WHEN "010110010101" => table_out <= 3576;
			WHEN "010110010110" => table_out <= 3577;
			WHEN "010110010111" => table_out <= 3577;
			WHEN "010110011000" => table_out <= 3577;
			WHEN "010110011001" => table_out <= 3578;
			WHEN "010110011010" => table_out <= 3578;
			WHEN "010110011011" => table_out <= 3578;
			WHEN "010110011100" => table_out <= 3579;
			WHEN "010110011101" => table_out <= 3579;
			WHEN "010110011110" => table_out <= 3579;
			WHEN "010110011111" => table_out <= 3580;
			WHEN "010110100000" => table_out <= 3580;
			WHEN "010110100001" => table_out <= 3580;
			WHEN "010110100010" => table_out <= 3581;
			WHEN "010110100011" => table_out <= 3581;
			WHEN "010110100100" => table_out <= 3581;
			WHEN "010110100101" => table_out <= 3582;
			WHEN "010110100110" => table_out <= 3582;
			WHEN "010110100111" => table_out <= 3582;
			WHEN "010110101000" => table_out <= 3583;
			WHEN "010110101001" => table_out <= 3583;
			WHEN "010110101010" => table_out <= 3583;
			WHEN "010110101011" => table_out <= 3584;
			WHEN "010110101100" => table_out <= 3584;
			WHEN "010110101101" => table_out <= 3584;
			WHEN "010110101110" => table_out <= 3585;
			WHEN "010110101111" => table_out <= 3585;
			WHEN "010110110000" => table_out <= 3586;
			WHEN "010110110001" => table_out <= 3586;
			WHEN "010110110010" => table_out <= 3586;
			WHEN "010110110011" => table_out <= 3587;
			WHEN "010110110100" => table_out <= 3587;
			WHEN "010110110101" => table_out <= 3587;
			WHEN "010110110110" => table_out <= 3588;
			WHEN "010110110111" => table_out <= 3588;
			WHEN "010110111000" => table_out <= 3588;
			WHEN "010110111001" => table_out <= 3589;
			WHEN "010110111010" => table_out <= 3589;
			WHEN "010110111011" => table_out <= 3589;
			WHEN "010110111100" => table_out <= 3590;
			WHEN "010110111101" => table_out <= 3590;
			WHEN "010110111110" => table_out <= 3590;
			WHEN "010110111111" => table_out <= 3591;
			WHEN "010111000000" => table_out <= 3591;
			WHEN "010111000001" => table_out <= 3591;
			WHEN "010111000010" => table_out <= 3592;
			WHEN "010111000011" => table_out <= 3592;
			WHEN "010111000100" => table_out <= 3592;
			WHEN "010111000101" => table_out <= 3593;
			WHEN "010111000110" => table_out <= 3593;
			WHEN "010111000111" => table_out <= 3593;
			WHEN "010111001000" => table_out <= 3594;
			WHEN "010111001001" => table_out <= 3594;
			WHEN "010111001010" => table_out <= 3594;
			WHEN "010111001011" => table_out <= 3595;
			WHEN "010111001100" => table_out <= 3595;
			WHEN "010111001101" => table_out <= 3595;
			WHEN "010111001110" => table_out <= 3596;
			WHEN "010111001111" => table_out <= 3596;
			WHEN "010111010000" => table_out <= 3596;
			WHEN "010111010001" => table_out <= 3597;
			WHEN "010111010010" => table_out <= 3597;
			WHEN "010111010011" => table_out <= 3597;
			WHEN "010111010100" => table_out <= 3598;
			WHEN "010111010101" => table_out <= 3598;
			WHEN "010111010110" => table_out <= 3598;
			WHEN "010111010111" => table_out <= 3599;
			WHEN "010111011000" => table_out <= 3599;
			WHEN "010111011001" => table_out <= 3599;
			WHEN "010111011010" => table_out <= 3600;
			WHEN "010111011011" => table_out <= 3600;
			WHEN "010111011100" => table_out <= 3600;
			WHEN "010111011101" => table_out <= 3600;
			WHEN "010111011110" => table_out <= 3601;
			WHEN "010111011111" => table_out <= 3601;
			WHEN "010111100000" => table_out <= 3601;
			WHEN "010111100001" => table_out <= 3602;
			WHEN "010111100010" => table_out <= 3602;
			WHEN "010111100011" => table_out <= 3602;
			WHEN "010111100100" => table_out <= 3603;
			WHEN "010111100101" => table_out <= 3603;
			WHEN "010111100110" => table_out <= 3603;
			WHEN "010111100111" => table_out <= 3604;
			WHEN "010111101000" => table_out <= 3604;
			WHEN "010111101001" => table_out <= 3604;
			WHEN "010111101010" => table_out <= 3605;
			WHEN "010111101011" => table_out <= 3605;
			WHEN "010111101100" => table_out <= 3605;
			WHEN "010111101101" => table_out <= 3606;
			WHEN "010111101110" => table_out <= 3606;
			WHEN "010111101111" => table_out <= 3606;
			WHEN "010111110000" => table_out <= 3607;
			WHEN "010111110001" => table_out <= 3607;
			WHEN "010111110010" => table_out <= 3607;
			WHEN "010111110011" => table_out <= 3608;
			WHEN "010111110100" => table_out <= 3608;
			WHEN "010111110101" => table_out <= 3608;
			WHEN "010111110110" => table_out <= 3609;
			WHEN "010111110111" => table_out <= 3609;
			WHEN "010111111000" => table_out <= 3609;
			WHEN "010111111001" => table_out <= 3610;
			WHEN "010111111010" => table_out <= 3610;
			WHEN "010111111011" => table_out <= 3610;
			WHEN "010111111100" => table_out <= 3611;
			WHEN "010111111101" => table_out <= 3611;
			WHEN "010111111110" => table_out <= 3611;
			WHEN "010111111111" => table_out <= 3612;
			WHEN "011000000000" => table_out <= 3612;
			WHEN "011000000001" => table_out <= 3612;
			WHEN "011000000010" => table_out <= 3612;
			WHEN "011000000011" => table_out <= 3613;
			WHEN "011000000100" => table_out <= 3613;
			WHEN "011000000101" => table_out <= 3613;
			WHEN "011000000110" => table_out <= 3614;
			WHEN "011000000111" => table_out <= 3614;
			WHEN "011000001000" => table_out <= 3614;
			WHEN "011000001001" => table_out <= 3615;
			WHEN "011000001010" => table_out <= 3615;
			WHEN "011000001011" => table_out <= 3615;
			WHEN "011000001100" => table_out <= 3616;
			WHEN "011000001101" => table_out <= 3616;
			WHEN "011000001110" => table_out <= 3616;
			WHEN "011000001111" => table_out <= 3617;
			WHEN "011000010000" => table_out <= 3617;
			WHEN "011000010001" => table_out <= 3617;
			WHEN "011000010010" => table_out <= 3618;
			WHEN "011000010011" => table_out <= 3618;
			WHEN "011000010100" => table_out <= 3618;
			WHEN "011000010101" => table_out <= 3619;
			WHEN "011000010110" => table_out <= 3619;
			WHEN "011000010111" => table_out <= 3619;
			WHEN "011000011000" => table_out <= 3619;
			WHEN "011000011001" => table_out <= 3620;
			WHEN "011000011010" => table_out <= 3620;
			WHEN "011000011011" => table_out <= 3620;
			WHEN "011000011100" => table_out <= 3621;
			WHEN "011000011101" => table_out <= 3621;
			WHEN "011000011110" => table_out <= 3621;
			WHEN "011000011111" => table_out <= 3622;
			WHEN "011000100000" => table_out <= 3622;
			WHEN "011000100001" => table_out <= 3622;
			WHEN "011000100010" => table_out <= 3623;
			WHEN "011000100011" => table_out <= 3623;
			WHEN "011000100100" => table_out <= 3623;
			WHEN "011000100101" => table_out <= 3624;
			WHEN "011000100110" => table_out <= 3624;
			WHEN "011000100111" => table_out <= 3624;
			WHEN "011000101000" => table_out <= 3624;
			WHEN "011000101001" => table_out <= 3625;
			WHEN "011000101010" => table_out <= 3625;
			WHEN "011000101011" => table_out <= 3625;
			WHEN "011000101100" => table_out <= 3626;
			WHEN "011000101101" => table_out <= 3626;
			WHEN "011000101110" => table_out <= 3626;
			WHEN "011000101111" => table_out <= 3627;
			WHEN "011000110000" => table_out <= 3627;
			WHEN "011000110001" => table_out <= 3627;
			WHEN "011000110010" => table_out <= 3628;
			WHEN "011000110011" => table_out <= 3628;
			WHEN "011000110100" => table_out <= 3628;
			WHEN "011000110101" => table_out <= 3629;
			WHEN "011000110110" => table_out <= 3629;
			WHEN "011000110111" => table_out <= 3629;
			WHEN "011000111000" => table_out <= 3629;
			WHEN "011000111001" => table_out <= 3630;
			WHEN "011000111010" => table_out <= 3630;
			WHEN "011000111011" => table_out <= 3630;
			WHEN "011000111100" => table_out <= 3631;
			WHEN "011000111101" => table_out <= 3631;
			WHEN "011000111110" => table_out <= 3631;
			WHEN "011000111111" => table_out <= 3632;
			WHEN "011001000000" => table_out <= 3632;
			WHEN "011001000001" => table_out <= 3632;
			WHEN "011001000010" => table_out <= 3633;
			WHEN "011001000011" => table_out <= 3633;
			WHEN "011001000100" => table_out <= 3633;
			WHEN "011001000101" => table_out <= 3633;
			WHEN "011001000110" => table_out <= 3634;
			WHEN "011001000111" => table_out <= 3634;
			WHEN "011001001000" => table_out <= 3634;
			WHEN "011001001001" => table_out <= 3635;
			WHEN "011001001010" => table_out <= 3635;
			WHEN "011001001011" => table_out <= 3635;
			WHEN "011001001100" => table_out <= 3636;
			WHEN "011001001101" => table_out <= 3636;
			WHEN "011001001110" => table_out <= 3636;
			WHEN "011001001111" => table_out <= 3637;
			WHEN "011001010000" => table_out <= 3637;
			WHEN "011001010001" => table_out <= 3637;
			WHEN "011001010010" => table_out <= 3637;
			WHEN "011001010011" => table_out <= 3638;
			WHEN "011001010100" => table_out <= 3638;
			WHEN "011001010101" => table_out <= 3638;
			WHEN "011001010110" => table_out <= 3639;
			WHEN "011001010111" => table_out <= 3639;
			WHEN "011001011000" => table_out <= 3639;
			WHEN "011001011001" => table_out <= 3640;
			WHEN "011001011010" => table_out <= 3640;
			WHEN "011001011011" => table_out <= 3640;
			WHEN "011001011100" => table_out <= 3640;
			WHEN "011001011101" => table_out <= 3641;
			WHEN "011001011110" => table_out <= 3641;
			WHEN "011001011111" => table_out <= 3641;
			WHEN "011001100000" => table_out <= 3642;
			WHEN "011001100001" => table_out <= 3642;
			WHEN "011001100010" => table_out <= 3642;
			WHEN "011001100011" => table_out <= 3643;
			WHEN "011001100100" => table_out <= 3643;
			WHEN "011001100101" => table_out <= 3643;
			WHEN "011001100110" => table_out <= 3643;
			WHEN "011001100111" => table_out <= 3644;
			WHEN "011001101000" => table_out <= 3644;
			WHEN "011001101001" => table_out <= 3644;
			WHEN "011001101010" => table_out <= 3645;
			WHEN "011001101011" => table_out <= 3645;
			WHEN "011001101100" => table_out <= 3645;
			WHEN "011001101101" => table_out <= 3646;
			WHEN "011001101110" => table_out <= 3646;
			WHEN "011001101111" => table_out <= 3646;
			WHEN "011001110000" => table_out <= 3646;
			WHEN "011001110001" => table_out <= 3647;
			WHEN "011001110010" => table_out <= 3647;
			WHEN "011001110011" => table_out <= 3647;
			WHEN "011001110100" => table_out <= 3648;
			WHEN "011001110101" => table_out <= 3648;
			WHEN "011001110110" => table_out <= 3648;
			WHEN "011001110111" => table_out <= 3649;
			WHEN "011001111000" => table_out <= 3649;
			WHEN "011001111001" => table_out <= 3649;
			WHEN "011001111010" => table_out <= 3649;
			WHEN "011001111011" => table_out <= 3650;
			WHEN "011001111100" => table_out <= 3650;
			WHEN "011001111101" => table_out <= 3650;
			WHEN "011001111110" => table_out <= 3651;
			WHEN "011001111111" => table_out <= 3651;
			WHEN "011010000000" => table_out <= 3651;
			WHEN "011010000001" => table_out <= 3652;
			WHEN "011010000010" => table_out <= 3652;
			WHEN "011010000011" => table_out <= 3652;
			WHEN "011010000100" => table_out <= 3652;
			WHEN "011010000101" => table_out <= 3653;
			WHEN "011010000110" => table_out <= 3653;
			WHEN "011010000111" => table_out <= 3653;
			WHEN "011010001000" => table_out <= 3654;
			WHEN "011010001001" => table_out <= 3654;
			WHEN "011010001010" => table_out <= 3654;
			WHEN "011010001011" => table_out <= 3654;
			WHEN "011010001100" => table_out <= 3655;
			WHEN "011010001101" => table_out <= 3655;
			WHEN "011010001110" => table_out <= 3655;
			WHEN "011010001111" => table_out <= 3656;
			WHEN "011010010000" => table_out <= 3656;
			WHEN "011010010001" => table_out <= 3656;
			WHEN "011010010010" => table_out <= 3657;
			WHEN "011010010011" => table_out <= 3657;
			WHEN "011010010100" => table_out <= 3657;
			WHEN "011010010101" => table_out <= 3657;
			WHEN "011010010110" => table_out <= 3658;
			WHEN "011010010111" => table_out <= 3658;
			WHEN "011010011000" => table_out <= 3658;
			WHEN "011010011001" => table_out <= 3659;
			WHEN "011010011010" => table_out <= 3659;
			WHEN "011010011011" => table_out <= 3659;
			WHEN "011010011100" => table_out <= 3659;
			WHEN "011010011101" => table_out <= 3660;
			WHEN "011010011110" => table_out <= 3660;
			WHEN "011010011111" => table_out <= 3660;
			WHEN "011010100000" => table_out <= 3661;
			WHEN "011010100001" => table_out <= 3661;
			WHEN "011010100010" => table_out <= 3661;
			WHEN "011010100011" => table_out <= 3661;
			WHEN "011010100100" => table_out <= 3662;
			WHEN "011010100101" => table_out <= 3662;
			WHEN "011010100110" => table_out <= 3662;
			WHEN "011010100111" => table_out <= 3663;
			WHEN "011010101000" => table_out <= 3663;
			WHEN "011010101001" => table_out <= 3663;
			WHEN "011010101010" => table_out <= 3664;
			WHEN "011010101011" => table_out <= 3664;
			WHEN "011010101100" => table_out <= 3664;
			WHEN "011010101101" => table_out <= 3664;
			WHEN "011010101110" => table_out <= 3665;
			WHEN "011010101111" => table_out <= 3665;
			WHEN "011010110000" => table_out <= 3665;
			WHEN "011010110001" => table_out <= 3666;
			WHEN "011010110010" => table_out <= 3666;
			WHEN "011010110011" => table_out <= 3666;
			WHEN "011010110100" => table_out <= 3666;
			WHEN "011010110101" => table_out <= 3667;
			WHEN "011010110110" => table_out <= 3667;
			WHEN "011010110111" => table_out <= 3667;
			WHEN "011010111000" => table_out <= 3668;
			WHEN "011010111001" => table_out <= 3668;
			WHEN "011010111010" => table_out <= 3668;
			WHEN "011010111011" => table_out <= 3668;
			WHEN "011010111100" => table_out <= 3669;
			WHEN "011010111101" => table_out <= 3669;
			WHEN "011010111110" => table_out <= 3669;
			WHEN "011010111111" => table_out <= 3670;
			WHEN "011011000000" => table_out <= 3670;
			WHEN "011011000001" => table_out <= 3670;
			WHEN "011011000010" => table_out <= 3670;
			WHEN "011011000011" => table_out <= 3671;
			WHEN "011011000100" => table_out <= 3671;
			WHEN "011011000101" => table_out <= 3671;
			WHEN "011011000110" => table_out <= 3672;
			WHEN "011011000111" => table_out <= 3672;
			WHEN "011011001000" => table_out <= 3672;
			WHEN "011011001001" => table_out <= 3672;
			WHEN "011011001010" => table_out <= 3673;
			WHEN "011011001011" => table_out <= 3673;
			WHEN "011011001100" => table_out <= 3673;
			WHEN "011011001101" => table_out <= 3674;
			WHEN "011011001110" => table_out <= 3674;
			WHEN "011011001111" => table_out <= 3674;
			WHEN "011011010000" => table_out <= 3674;
			WHEN "011011010001" => table_out <= 3675;
			WHEN "011011010010" => table_out <= 3675;
			WHEN "011011010011" => table_out <= 3675;
			WHEN "011011010100" => table_out <= 3675;
			WHEN "011011010101" => table_out <= 3676;
			WHEN "011011010110" => table_out <= 3676;
			WHEN "011011010111" => table_out <= 3676;
			WHEN "011011011000" => table_out <= 3677;
			WHEN "011011011001" => table_out <= 3677;
			WHEN "011011011010" => table_out <= 3677;
			WHEN "011011011011" => table_out <= 3677;
			WHEN "011011011100" => table_out <= 3678;
			WHEN "011011011101" => table_out <= 3678;
			WHEN "011011011110" => table_out <= 3678;
			WHEN "011011011111" => table_out <= 3679;
			WHEN "011011100000" => table_out <= 3679;
			WHEN "011011100001" => table_out <= 3679;
			WHEN "011011100010" => table_out <= 3679;
			WHEN "011011100011" => table_out <= 3680;
			WHEN "011011100100" => table_out <= 3680;
			WHEN "011011100101" => table_out <= 3680;
			WHEN "011011100110" => table_out <= 3681;
			WHEN "011011100111" => table_out <= 3681;
			WHEN "011011101000" => table_out <= 3681;
			WHEN "011011101001" => table_out <= 3681;
			WHEN "011011101010" => table_out <= 3682;
			WHEN "011011101011" => table_out <= 3682;
			WHEN "011011101100" => table_out <= 3682;
			WHEN "011011101101" => table_out <= 3682;
			WHEN "011011101110" => table_out <= 3683;
			WHEN "011011101111" => table_out <= 3683;
			WHEN "011011110000" => table_out <= 3683;
			WHEN "011011110001" => table_out <= 3684;
			WHEN "011011110010" => table_out <= 3684;
			WHEN "011011110011" => table_out <= 3684;
			WHEN "011011110100" => table_out <= 3684;
			WHEN "011011110101" => table_out <= 3685;
			WHEN "011011110110" => table_out <= 3685;
			WHEN "011011110111" => table_out <= 3685;
			WHEN "011011111000" => table_out <= 3686;
			WHEN "011011111001" => table_out <= 3686;
			WHEN "011011111010" => table_out <= 3686;
			WHEN "011011111011" => table_out <= 3686;
			WHEN "011011111100" => table_out <= 3687;
			WHEN "011011111101" => table_out <= 3687;
			WHEN "011011111110" => table_out <= 3687;
			WHEN "011011111111" => table_out <= 3687;
			WHEN "011100000000" => table_out <= 3688;
			WHEN "011100000001" => table_out <= 3688;
			WHEN "011100000010" => table_out <= 3688;
			WHEN "011100000011" => table_out <= 3689;
			WHEN "011100000100" => table_out <= 3689;
			WHEN "011100000101" => table_out <= 3689;
			WHEN "011100000110" => table_out <= 3689;
			WHEN "011100000111" => table_out <= 3690;
			WHEN "011100001000" => table_out <= 3690;
			WHEN "011100001001" => table_out <= 3690;
			WHEN "011100001010" => table_out <= 3690;
			WHEN "011100001011" => table_out <= 3691;
			WHEN "011100001100" => table_out <= 3691;
			WHEN "011100001101" => table_out <= 3691;
			WHEN "011100001110" => table_out <= 3692;
			WHEN "011100001111" => table_out <= 3692;
			WHEN "011100010000" => table_out <= 3692;
			WHEN "011100010001" => table_out <= 3692;
			WHEN "011100010010" => table_out <= 3693;
			WHEN "011100010011" => table_out <= 3693;
			WHEN "011100010100" => table_out <= 3693;
			WHEN "011100010101" => table_out <= 3693;
			WHEN "011100010110" => table_out <= 3694;
			WHEN "011100010111" => table_out <= 3694;
			WHEN "011100011000" => table_out <= 3694;
			WHEN "011100011001" => table_out <= 3695;
			WHEN "011100011010" => table_out <= 3695;
			WHEN "011100011011" => table_out <= 3695;
			WHEN "011100011100" => table_out <= 3695;
			WHEN "011100011101" => table_out <= 3696;
			WHEN "011100011110" => table_out <= 3696;
			WHEN "011100011111" => table_out <= 3696;
			WHEN "011100100000" => table_out <= 3696;
			WHEN "011100100001" => table_out <= 3697;
			WHEN "011100100010" => table_out <= 3697;
			WHEN "011100100011" => table_out <= 3697;
			WHEN "011100100100" => table_out <= 3698;
			WHEN "011100100101" => table_out <= 3698;
			WHEN "011100100110" => table_out <= 3698;
			WHEN "011100100111" => table_out <= 3698;
			WHEN "011100101000" => table_out <= 3699;
			WHEN "011100101001" => table_out <= 3699;
			WHEN "011100101010" => table_out <= 3699;
			WHEN "011100101011" => table_out <= 3699;
			WHEN "011100101100" => table_out <= 3700;
			WHEN "011100101101" => table_out <= 3700;
			WHEN "011100101110" => table_out <= 3700;
			WHEN "011100101111" => table_out <= 3700;
			WHEN "011100110000" => table_out <= 3701;
			WHEN "011100110001" => table_out <= 3701;
			WHEN "011100110010" => table_out <= 3701;
			WHEN "011100110011" => table_out <= 3702;
			WHEN "011100110100" => table_out <= 3702;
			WHEN "011100110101" => table_out <= 3702;
			WHEN "011100110110" => table_out <= 3702;
			WHEN "011100110111" => table_out <= 3703;
			WHEN "011100111000" => table_out <= 3703;
			WHEN "011100111001" => table_out <= 3703;
			WHEN "011100111010" => table_out <= 3703;
			WHEN "011100111011" => table_out <= 3704;
			WHEN "011100111100" => table_out <= 3704;
			WHEN "011100111101" => table_out <= 3704;
			WHEN "011100111110" => table_out <= 3704;
			WHEN "011100111111" => table_out <= 3705;
			WHEN "011101000000" => table_out <= 3705;
			WHEN "011101000001" => table_out <= 3705;
			WHEN "011101000010" => table_out <= 3706;
			WHEN "011101000011" => table_out <= 3706;
			WHEN "011101000100" => table_out <= 3706;
			WHEN "011101000101" => table_out <= 3706;
			WHEN "011101000110" => table_out <= 3707;
			WHEN "011101000111" => table_out <= 3707;
			WHEN "011101001000" => table_out <= 3707;
			WHEN "011101001001" => table_out <= 3707;
			WHEN "011101001010" => table_out <= 3708;
			WHEN "011101001011" => table_out <= 3708;
			WHEN "011101001100" => table_out <= 3708;
			WHEN "011101001101" => table_out <= 3708;
			WHEN "011101001110" => table_out <= 3709;
			WHEN "011101001111" => table_out <= 3709;
			WHEN "011101010000" => table_out <= 3709;
			WHEN "011101010001" => table_out <= 3709;
			WHEN "011101010010" => table_out <= 3710;
			WHEN "011101010011" => table_out <= 3710;
			WHEN "011101010100" => table_out <= 3710;
			WHEN "011101010101" => table_out <= 3711;
			WHEN "011101010110" => table_out <= 3711;
			WHEN "011101010111" => table_out <= 3711;
			WHEN "011101011000" => table_out <= 3711;
			WHEN "011101011001" => table_out <= 3712;
			WHEN "011101011010" => table_out <= 3712;
			WHEN "011101011011" => table_out <= 3712;
			WHEN "011101011100" => table_out <= 3712;
			WHEN "011101011101" => table_out <= 3713;
			WHEN "011101011110" => table_out <= 3713;
			WHEN "011101011111" => table_out <= 3713;
			WHEN "011101100000" => table_out <= 3713;
			WHEN "011101100001" => table_out <= 3714;
			WHEN "011101100010" => table_out <= 3714;
			WHEN "011101100011" => table_out <= 3714;
			WHEN "011101100100" => table_out <= 3714;
			WHEN "011101100101" => table_out <= 3715;
			WHEN "011101100110" => table_out <= 3715;
			WHEN "011101100111" => table_out <= 3715;
			WHEN "011101101000" => table_out <= 3715;
			WHEN "011101101001" => table_out <= 3716;
			WHEN "011101101010" => table_out <= 3716;
			WHEN "011101101011" => table_out <= 3716;
			WHEN "011101101100" => table_out <= 3717;
			WHEN "011101101101" => table_out <= 3717;
			WHEN "011101101110" => table_out <= 3717;
			WHEN "011101101111" => table_out <= 3717;
			WHEN "011101110000" => table_out <= 3718;
			WHEN "011101110001" => table_out <= 3718;
			WHEN "011101110010" => table_out <= 3718;
			WHEN "011101110011" => table_out <= 3718;
			WHEN "011101110100" => table_out <= 3719;
			WHEN "011101110101" => table_out <= 3719;
			WHEN "011101110110" => table_out <= 3719;
			WHEN "011101110111" => table_out <= 3719;
			WHEN "011101111000" => table_out <= 3720;
			WHEN "011101111001" => table_out <= 3720;
			WHEN "011101111010" => table_out <= 3720;
			WHEN "011101111011" => table_out <= 3720;
			WHEN "011101111100" => table_out <= 3721;
			WHEN "011101111101" => table_out <= 3721;
			WHEN "011101111110" => table_out <= 3721;
			WHEN "011101111111" => table_out <= 3721;
			WHEN "011110000000" => table_out <= 3722;
			WHEN "011110000001" => table_out <= 3722;
			WHEN "011110000010" => table_out <= 3722;
			WHEN "011110000011" => table_out <= 3722;
			WHEN "011110000100" => table_out <= 3723;
			WHEN "011110000101" => table_out <= 3723;
			WHEN "011110000110" => table_out <= 3723;
			WHEN "011110000111" => table_out <= 3723;
			WHEN "011110001000" => table_out <= 3724;
			WHEN "011110001001" => table_out <= 3724;
			WHEN "011110001010" => table_out <= 3724;
			WHEN "011110001011" => table_out <= 3724;
			WHEN "011110001100" => table_out <= 3725;
			WHEN "011110001101" => table_out <= 3725;
			WHEN "011110001110" => table_out <= 3725;
			WHEN "011110001111" => table_out <= 3726;
			WHEN "011110010000" => table_out <= 3726;
			WHEN "011110010001" => table_out <= 3726;
			WHEN "011110010010" => table_out <= 3726;
			WHEN "011110010011" => table_out <= 3727;
			WHEN "011110010100" => table_out <= 3727;
			WHEN "011110010101" => table_out <= 3727;
			WHEN "011110010110" => table_out <= 3727;
			WHEN "011110010111" => table_out <= 3728;
			WHEN "011110011000" => table_out <= 3728;
			WHEN "011110011001" => table_out <= 3728;
			WHEN "011110011010" => table_out <= 3728;
			WHEN "011110011011" => table_out <= 3729;
			WHEN "011110011100" => table_out <= 3729;
			WHEN "011110011101" => table_out <= 3729;
			WHEN "011110011110" => table_out <= 3729;
			WHEN "011110011111" => table_out <= 3730;
			WHEN "011110100000" => table_out <= 3730;
			WHEN "011110100001" => table_out <= 3730;
			WHEN "011110100010" => table_out <= 3730;
			WHEN "011110100011" => table_out <= 3731;
			WHEN "011110100100" => table_out <= 3731;
			WHEN "011110100101" => table_out <= 3731;
			WHEN "011110100110" => table_out <= 3731;
			WHEN "011110100111" => table_out <= 3732;
			WHEN "011110101000" => table_out <= 3732;
			WHEN "011110101001" => table_out <= 3732;
			WHEN "011110101010" => table_out <= 3732;
			WHEN "011110101011" => table_out <= 3733;
			WHEN "011110101100" => table_out <= 3733;
			WHEN "011110101101" => table_out <= 3733;
			WHEN "011110101110" => table_out <= 3733;
			WHEN "011110101111" => table_out <= 3734;
			WHEN "011110110000" => table_out <= 3734;
			WHEN "011110110001" => table_out <= 3734;
			WHEN "011110110010" => table_out <= 3734;
			WHEN "011110110011" => table_out <= 3735;
			WHEN "011110110100" => table_out <= 3735;
			WHEN "011110110101" => table_out <= 3735;
			WHEN "011110110110" => table_out <= 3735;
			WHEN "011110110111" => table_out <= 3736;
			WHEN "011110111000" => table_out <= 3736;
			WHEN "011110111001" => table_out <= 3736;
			WHEN "011110111010" => table_out <= 3736;
			WHEN "011110111011" => table_out <= 3737;
			WHEN "011110111100" => table_out <= 3737;
			WHEN "011110111101" => table_out <= 3737;
			WHEN "011110111110" => table_out <= 3737;
			WHEN "011110111111" => table_out <= 3738;
			WHEN "011111000000" => table_out <= 3738;
			WHEN "011111000001" => table_out <= 3738;
			WHEN "011111000010" => table_out <= 3738;
			WHEN "011111000011" => table_out <= 3739;
			WHEN "011111000100" => table_out <= 3739;
			WHEN "011111000101" => table_out <= 3739;
			WHEN "011111000110" => table_out <= 3739;
			WHEN "011111000111" => table_out <= 3740;
			WHEN "011111001000" => table_out <= 3740;
			WHEN "011111001001" => table_out <= 3740;
			WHEN "011111001010" => table_out <= 3740;
			WHEN "011111001011" => table_out <= 3741;
			WHEN "011111001100" => table_out <= 3741;
			WHEN "011111001101" => table_out <= 3741;
			WHEN "011111001110" => table_out <= 3741;
			WHEN "011111001111" => table_out <= 3742;
			WHEN "011111010000" => table_out <= 3742;
			WHEN "011111010001" => table_out <= 3742;
			WHEN "011111010010" => table_out <= 3742;
			WHEN "011111010011" => table_out <= 3743;
			WHEN "011111010100" => table_out <= 3743;
			WHEN "011111010101" => table_out <= 3743;
			WHEN "011111010110" => table_out <= 3743;
			WHEN "011111010111" => table_out <= 3743;
			WHEN "011111011000" => table_out <= 3744;
			WHEN "011111011001" => table_out <= 3744;
			WHEN "011111011010" => table_out <= 3744;
			WHEN "011111011011" => table_out <= 3744;
			WHEN "011111011100" => table_out <= 3745;
			WHEN "011111011101" => table_out <= 3745;
			WHEN "011111011110" => table_out <= 3745;
			WHEN "011111011111" => table_out <= 3745;
			WHEN "011111100000" => table_out <= 3746;
			WHEN "011111100001" => table_out <= 3746;
			WHEN "011111100010" => table_out <= 3746;
			WHEN "011111100011" => table_out <= 3746;
			WHEN "011111100100" => table_out <= 3747;
			WHEN "011111100101" => table_out <= 3747;
			WHEN "011111100110" => table_out <= 3747;
			WHEN "011111100111" => table_out <= 3747;
			WHEN "011111101000" => table_out <= 3748;
			WHEN "011111101001" => table_out <= 3748;
			WHEN "011111101010" => table_out <= 3748;
			WHEN "011111101011" => table_out <= 3748;
			WHEN "011111101100" => table_out <= 3749;
			WHEN "011111101101" => table_out <= 3749;
			WHEN "011111101110" => table_out <= 3749;
			WHEN "011111101111" => table_out <= 3749;
			WHEN "011111110000" => table_out <= 3750;
			WHEN "011111110001" => table_out <= 3750;
			WHEN "011111110010" => table_out <= 3750;
			WHEN "011111110011" => table_out <= 3750;
			WHEN "011111110100" => table_out <= 3751;
			WHEN "011111110101" => table_out <= 3751;
			WHEN "011111110110" => table_out <= 3751;
			WHEN "011111110111" => table_out <= 3751;
			WHEN "011111111000" => table_out <= 3752;
			WHEN "011111111001" => table_out <= 3752;
			WHEN "011111111010" => table_out <= 3752;
			WHEN "011111111011" => table_out <= 3752;
			WHEN "011111111100" => table_out <= 3752;
			WHEN "011111111101" => table_out <= 3753;
			WHEN "011111111110" => table_out <= 3753;
			WHEN "011111111111" => table_out <= 3753;
			WHEN "100000000000" => table_out <= 3753;
			WHEN "100000000001" => table_out <= 3754;
			WHEN "100000000010" => table_out <= 3754;
			WHEN "100000000011" => table_out <= 3754;
			WHEN "100000000100" => table_out <= 3754;
			WHEN "100000000101" => table_out <= 3755;
			WHEN "100000000110" => table_out <= 3755;
			WHEN "100000000111" => table_out <= 3755;
			WHEN "100000001000" => table_out <= 3755;
			WHEN "100000001001" => table_out <= 3756;
			WHEN "100000001010" => table_out <= 3756;
			WHEN "100000001011" => table_out <= 3756;
			WHEN "100000001100" => table_out <= 3756;
			WHEN "100000001101" => table_out <= 3757;
			WHEN "100000001110" => table_out <= 3757;
			WHEN "100000001111" => table_out <= 3757;
			WHEN "100000010000" => table_out <= 3757;
			WHEN "100000010001" => table_out <= 3758;
			WHEN "100000010010" => table_out <= 3758;
			WHEN "100000010011" => table_out <= 3758;
			WHEN "100000010100" => table_out <= 3758;
			WHEN "100000010101" => table_out <= 3758;
			WHEN "100000010110" => table_out <= 3759;
			WHEN "100000010111" => table_out <= 3759;
			WHEN "100000011000" => table_out <= 3759;
			WHEN "100000011001" => table_out <= 3759;
			WHEN "100000011010" => table_out <= 3760;
			WHEN "100000011011" => table_out <= 3760;
			WHEN "100000011100" => table_out <= 3760;
			WHEN "100000011101" => table_out <= 3760;
			WHEN "100000011110" => table_out <= 3761;
			WHEN "100000011111" => table_out <= 3761;
			WHEN "100000100000" => table_out <= 3761;
			WHEN "100000100001" => table_out <= 3761;
			WHEN "100000100010" => table_out <= 3762;
			WHEN "100000100011" => table_out <= 3762;
			WHEN "100000100100" => table_out <= 3762;
			WHEN "100000100101" => table_out <= 3762;
			WHEN "100000100110" => table_out <= 3762;
			WHEN "100000100111" => table_out <= 3763;
			WHEN "100000101000" => table_out <= 3763;
			WHEN "100000101001" => table_out <= 3763;
			WHEN "100000101010" => table_out <= 3763;
			WHEN "100000101011" => table_out <= 3764;
			WHEN "100000101100" => table_out <= 3764;
			WHEN "100000101101" => table_out <= 3764;
			WHEN "100000101110" => table_out <= 3764;
			WHEN "100000101111" => table_out <= 3765;
			WHEN "100000110000" => table_out <= 3765;
			WHEN "100000110001" => table_out <= 3765;
			WHEN "100000110010" => table_out <= 3765;
			WHEN "100000110011" => table_out <= 3766;
			WHEN "100000110100" => table_out <= 3766;
			WHEN "100000110101" => table_out <= 3766;
			WHEN "100000110110" => table_out <= 3766;
			WHEN "100000110111" => table_out <= 3766;
			WHEN "100000111000" => table_out <= 3767;
			WHEN "100000111001" => table_out <= 3767;
			WHEN "100000111010" => table_out <= 3767;
			WHEN "100000111011" => table_out <= 3767;
			WHEN "100000111100" => table_out <= 3768;
			WHEN "100000111101" => table_out <= 3768;
			WHEN "100000111110" => table_out <= 3768;
			WHEN "100000111111" => table_out <= 3768;
			WHEN "100001000000" => table_out <= 3769;
			WHEN "100001000001" => table_out <= 3769;
			WHEN "100001000010" => table_out <= 3769;
			WHEN "100001000011" => table_out <= 3769;
			WHEN "100001000100" => table_out <= 3770;
			WHEN "100001000101" => table_out <= 3770;
			WHEN "100001000110" => table_out <= 3770;
			WHEN "100001000111" => table_out <= 3770;
			WHEN "100001001000" => table_out <= 3770;
			WHEN "100001001001" => table_out <= 3771;
			WHEN "100001001010" => table_out <= 3771;
			WHEN "100001001011" => table_out <= 3771;
			WHEN "100001001100" => table_out <= 3771;
			WHEN "100001001101" => table_out <= 3772;
			WHEN "100001001110" => table_out <= 3772;
			WHEN "100001001111" => table_out <= 3772;
			WHEN "100001010000" => table_out <= 3772;
			WHEN "100001010001" => table_out <= 3773;
			WHEN "100001010010" => table_out <= 3773;
			WHEN "100001010011" => table_out <= 3773;
			WHEN "100001010100" => table_out <= 3773;
			WHEN "100001010101" => table_out <= 3773;
			WHEN "100001010110" => table_out <= 3774;
			WHEN "100001010111" => table_out <= 3774;
			WHEN "100001011000" => table_out <= 3774;
			WHEN "100001011001" => table_out <= 3774;
			WHEN "100001011010" => table_out <= 3775;
			WHEN "100001011011" => table_out <= 3775;
			WHEN "100001011100" => table_out <= 3775;
			WHEN "100001011101" => table_out <= 3775;
			WHEN "100001011110" => table_out <= 3776;
			WHEN "100001011111" => table_out <= 3776;
			WHEN "100001100000" => table_out <= 3776;
			WHEN "100001100001" => table_out <= 3776;
			WHEN "100001100010" => table_out <= 3776;
			WHEN "100001100011" => table_out <= 3777;
			WHEN "100001100100" => table_out <= 3777;
			WHEN "100001100101" => table_out <= 3777;
			WHEN "100001100110" => table_out <= 3777;
			WHEN "100001100111" => table_out <= 3778;
			WHEN "100001101000" => table_out <= 3778;
			WHEN "100001101001" => table_out <= 3778;
			WHEN "100001101010" => table_out <= 3778;
			WHEN "100001101011" => table_out <= 3779;
			WHEN "100001101100" => table_out <= 3779;
			WHEN "100001101101" => table_out <= 3779;
			WHEN "100001101110" => table_out <= 3779;
			WHEN "100001101111" => table_out <= 3779;
			WHEN "100001110000" => table_out <= 3780;
			WHEN "100001110001" => table_out <= 3780;
			WHEN "100001110010" => table_out <= 3780;
			WHEN "100001110011" => table_out <= 3780;
			WHEN "100001110100" => table_out <= 3781;
			WHEN "100001110101" => table_out <= 3781;
			WHEN "100001110110" => table_out <= 3781;
			WHEN "100001110111" => table_out <= 3781;
			WHEN "100001111000" => table_out <= 3781;
			WHEN "100001111001" => table_out <= 3782;
			WHEN "100001111010" => table_out <= 3782;
			WHEN "100001111011" => table_out <= 3782;
			WHEN "100001111100" => table_out <= 3782;
			WHEN "100001111101" => table_out <= 3783;
			WHEN "100001111110" => table_out <= 3783;
			WHEN "100001111111" => table_out <= 3783;
			WHEN "100010000000" => table_out <= 3783;
			WHEN "100010000001" => table_out <= 3784;
			WHEN "100010000010" => table_out <= 3784;
			WHEN "100010000011" => table_out <= 3784;
			WHEN "100010000100" => table_out <= 3784;
			WHEN "100010000101" => table_out <= 3784;
			WHEN "100010000110" => table_out <= 3785;
			WHEN "100010000111" => table_out <= 3785;
			WHEN "100010001000" => table_out <= 3785;
			WHEN "100010001001" => table_out <= 3785;
			WHEN "100010001010" => table_out <= 3786;
			WHEN "100010001011" => table_out <= 3786;
			WHEN "100010001100" => table_out <= 3786;
			WHEN "100010001101" => table_out <= 3786;
			WHEN "100010001110" => table_out <= 3786;
			WHEN "100010001111" => table_out <= 3787;
			WHEN "100010010000" => table_out <= 3787;
			WHEN "100010010001" => table_out <= 3787;
			WHEN "100010010010" => table_out <= 3787;
			WHEN "100010010011" => table_out <= 3788;
			WHEN "100010010100" => table_out <= 3788;
			WHEN "100010010101" => table_out <= 3788;
			WHEN "100010010110" => table_out <= 3788;
			WHEN "100010010111" => table_out <= 3788;
			WHEN "100010011000" => table_out <= 3789;
			WHEN "100010011001" => table_out <= 3789;
			WHEN "100010011010" => table_out <= 3789;
			WHEN "100010011011" => table_out <= 3789;
			WHEN "100010011100" => table_out <= 3790;
			WHEN "100010011101" => table_out <= 3790;
			WHEN "100010011110" => table_out <= 3790;
			WHEN "100010011111" => table_out <= 3790;
			WHEN "100010100000" => table_out <= 3790;
			WHEN "100010100001" => table_out <= 3791;
			WHEN "100010100010" => table_out <= 3791;
			WHEN "100010100011" => table_out <= 3791;
			WHEN "100010100100" => table_out <= 3791;
			WHEN "100010100101" => table_out <= 3792;
			WHEN "100010100110" => table_out <= 3792;
			WHEN "100010100111" => table_out <= 3792;
			WHEN "100010101000" => table_out <= 3792;
			WHEN "100010101001" => table_out <= 3792;
			WHEN "100010101010" => table_out <= 3793;
			WHEN "100010101011" => table_out <= 3793;
			WHEN "100010101100" => table_out <= 3793;
			WHEN "100010101101" => table_out <= 3793;
			WHEN "100010101110" => table_out <= 3794;
			WHEN "100010101111" => table_out <= 3794;
			WHEN "100010110000" => table_out <= 3794;
			WHEN "100010110001" => table_out <= 3794;
			WHEN "100010110010" => table_out <= 3794;
			WHEN "100010110011" => table_out <= 3795;
			WHEN "100010110100" => table_out <= 3795;
			WHEN "100010110101" => table_out <= 3795;
			WHEN "100010110110" => table_out <= 3795;
			WHEN "100010110111" => table_out <= 3796;
			WHEN "100010111000" => table_out <= 3796;
			WHEN "100010111001" => table_out <= 3796;
			WHEN "100010111010" => table_out <= 3796;
			WHEN "100010111011" => table_out <= 3796;
			WHEN "100010111100" => table_out <= 3797;
			WHEN "100010111101" => table_out <= 3797;
			WHEN "100010111110" => table_out <= 3797;
			WHEN "100010111111" => table_out <= 3797;
			WHEN "100011000000" => table_out <= 3798;
			WHEN "100011000001" => table_out <= 3798;
			WHEN "100011000010" => table_out <= 3798;
			WHEN "100011000011" => table_out <= 3798;
			WHEN "100011000100" => table_out <= 3798;
			WHEN "100011000101" => table_out <= 3799;
			WHEN "100011000110" => table_out <= 3799;
			WHEN "100011000111" => table_out <= 3799;
			WHEN "100011001000" => table_out <= 3799;
			WHEN "100011001001" => table_out <= 3800;
			WHEN "100011001010" => table_out <= 3800;
			WHEN "100011001011" => table_out <= 3800;
			WHEN "100011001100" => table_out <= 3800;
			WHEN "100011001101" => table_out <= 3800;
			WHEN "100011001110" => table_out <= 3801;
			WHEN "100011001111" => table_out <= 3801;
			WHEN "100011010000" => table_out <= 3801;
			WHEN "100011010001" => table_out <= 3801;
			WHEN "100011010010" => table_out <= 3801;
			WHEN "100011010011" => table_out <= 3802;
			WHEN "100011010100" => table_out <= 3802;
			WHEN "100011010101" => table_out <= 3802;
			WHEN "100011010110" => table_out <= 3802;
			WHEN "100011010111" => table_out <= 3803;
			WHEN "100011011000" => table_out <= 3803;
			WHEN "100011011001" => table_out <= 3803;
			WHEN "100011011010" => table_out <= 3803;
			WHEN "100011011011" => table_out <= 3803;
			WHEN "100011011100" => table_out <= 3804;
			WHEN "100011011101" => table_out <= 3804;
			WHEN "100011011110" => table_out <= 3804;
			WHEN "100011011111" => table_out <= 3804;
			WHEN "100011100000" => table_out <= 3805;
			WHEN "100011100001" => table_out <= 3805;
			WHEN "100011100010" => table_out <= 3805;
			WHEN "100011100011" => table_out <= 3805;
			WHEN "100011100100" => table_out <= 3805;
			WHEN "100011100101" => table_out <= 3806;
			WHEN "100011100110" => table_out <= 3806;
			WHEN "100011100111" => table_out <= 3806;
			WHEN "100011101000" => table_out <= 3806;
			WHEN "100011101001" => table_out <= 3806;
			WHEN "100011101010" => table_out <= 3807;
			WHEN "100011101011" => table_out <= 3807;
			WHEN "100011101100" => table_out <= 3807;
			WHEN "100011101101" => table_out <= 3807;
			WHEN "100011101110" => table_out <= 3808;
			WHEN "100011101111" => table_out <= 3808;
			WHEN "100011110000" => table_out <= 3808;
			WHEN "100011110001" => table_out <= 3808;
			WHEN "100011110010" => table_out <= 3808;
			WHEN "100011110011" => table_out <= 3809;
			WHEN "100011110100" => table_out <= 3809;
			WHEN "100011110101" => table_out <= 3809;
			WHEN "100011110110" => table_out <= 3809;
			WHEN "100011110111" => table_out <= 3809;
			WHEN "100011111000" => table_out <= 3810;
			WHEN "100011111001" => table_out <= 3810;
			WHEN "100011111010" => table_out <= 3810;
			WHEN "100011111011" => table_out <= 3810;
			WHEN "100011111100" => table_out <= 3811;
			WHEN "100011111101" => table_out <= 3811;
			WHEN "100011111110" => table_out <= 3811;
			WHEN "100011111111" => table_out <= 3811;
			WHEN "100100000000" => table_out <= 3811;
			WHEN "100100000001" => table_out <= 3812;
			WHEN "100100000010" => table_out <= 3812;
			WHEN "100100000011" => table_out <= 3812;
			WHEN "100100000100" => table_out <= 3812;
			WHEN "100100000101" => table_out <= 3812;
			WHEN "100100000110" => table_out <= 3813;
			WHEN "100100000111" => table_out <= 3813;
			WHEN "100100001000" => table_out <= 3813;
			WHEN "100100001001" => table_out <= 3813;
			WHEN "100100001010" => table_out <= 3814;
			WHEN "100100001011" => table_out <= 3814;
			WHEN "100100001100" => table_out <= 3814;
			WHEN "100100001101" => table_out <= 3814;
			WHEN "100100001110" => table_out <= 3814;
			WHEN "100100001111" => table_out <= 3815;
			WHEN "100100010000" => table_out <= 3815;
			WHEN "100100010001" => table_out <= 3815;
			WHEN "100100010010" => table_out <= 3815;
			WHEN "100100010011" => table_out <= 3815;
			WHEN "100100010100" => table_out <= 3816;
			WHEN "100100010101" => table_out <= 3816;
			WHEN "100100010110" => table_out <= 3816;
			WHEN "100100010111" => table_out <= 3816;
			WHEN "100100011000" => table_out <= 3817;
			WHEN "100100011001" => table_out <= 3817;
			WHEN "100100011010" => table_out <= 3817;
			WHEN "100100011011" => table_out <= 3817;
			WHEN "100100011100" => table_out <= 3817;
			WHEN "100100011101" => table_out <= 3818;
			WHEN "100100011110" => table_out <= 3818;
			WHEN "100100011111" => table_out <= 3818;
			WHEN "100100100000" => table_out <= 3818;
			WHEN "100100100001" => table_out <= 3818;
			WHEN "100100100010" => table_out <= 3819;
			WHEN "100100100011" => table_out <= 3819;
			WHEN "100100100100" => table_out <= 3819;
			WHEN "100100100101" => table_out <= 3819;
			WHEN "100100100110" => table_out <= 3819;
			WHEN "100100100111" => table_out <= 3820;
			WHEN "100100101000" => table_out <= 3820;
			WHEN "100100101001" => table_out <= 3820;
			WHEN "100100101010" => table_out <= 3820;
			WHEN "100100101011" => table_out <= 3821;
			WHEN "100100101100" => table_out <= 3821;
			WHEN "100100101101" => table_out <= 3821;
			WHEN "100100101110" => table_out <= 3821;
			WHEN "100100101111" => table_out <= 3821;
			WHEN "100100110000" => table_out <= 3822;
			WHEN "100100110001" => table_out <= 3822;
			WHEN "100100110010" => table_out <= 3822;
			WHEN "100100110011" => table_out <= 3822;
			WHEN "100100110100" => table_out <= 3822;
			WHEN "100100110101" => table_out <= 3823;
			WHEN "100100110110" => table_out <= 3823;
			WHEN "100100110111" => table_out <= 3823;
			WHEN "100100111000" => table_out <= 3823;
			WHEN "100100111001" => table_out <= 3823;
			WHEN "100100111010" => table_out <= 3824;
			WHEN "100100111011" => table_out <= 3824;
			WHEN "100100111100" => table_out <= 3824;
			WHEN "100100111101" => table_out <= 3824;
			WHEN "100100111110" => table_out <= 3824;
			WHEN "100100111111" => table_out <= 3825;
			WHEN "100101000000" => table_out <= 3825;
			WHEN "100101000001" => table_out <= 3825;
			WHEN "100101000010" => table_out <= 3825;
			WHEN "100101000011" => table_out <= 3826;
			WHEN "100101000100" => table_out <= 3826;
			WHEN "100101000101" => table_out <= 3826;
			WHEN "100101000110" => table_out <= 3826;
			WHEN "100101000111" => table_out <= 3826;
			WHEN "100101001000" => table_out <= 3827;
			WHEN "100101001001" => table_out <= 3827;
			WHEN "100101001010" => table_out <= 3827;
			WHEN "100101001011" => table_out <= 3827;
			WHEN "100101001100" => table_out <= 3827;
			WHEN "100101001101" => table_out <= 3828;
			WHEN "100101001110" => table_out <= 3828;
			WHEN "100101001111" => table_out <= 3828;
			WHEN "100101010000" => table_out <= 3828;
			WHEN "100101010001" => table_out <= 3828;
			WHEN "100101010010" => table_out <= 3829;
			WHEN "100101010011" => table_out <= 3829;
			WHEN "100101010100" => table_out <= 3829;
			WHEN "100101010101" => table_out <= 3829;
			WHEN "100101010110" => table_out <= 3829;
			WHEN "100101010111" => table_out <= 3830;
			WHEN "100101011000" => table_out <= 3830;
			WHEN "100101011001" => table_out <= 3830;
			WHEN "100101011010" => table_out <= 3830;
			WHEN "100101011011" => table_out <= 3830;
			WHEN "100101011100" => table_out <= 3831;
			WHEN "100101011101" => table_out <= 3831;
			WHEN "100101011110" => table_out <= 3831;
			WHEN "100101011111" => table_out <= 3831;
			WHEN "100101100000" => table_out <= 3832;
			WHEN "100101100001" => table_out <= 3832;
			WHEN "100101100010" => table_out <= 3832;
			WHEN "100101100011" => table_out <= 3832;
			WHEN "100101100100" => table_out <= 3832;
			WHEN "100101100101" => table_out <= 3833;
			WHEN "100101100110" => table_out <= 3833;
			WHEN "100101100111" => table_out <= 3833;
			WHEN "100101101000" => table_out <= 3833;
			WHEN "100101101001" => table_out <= 3833;
			WHEN "100101101010" => table_out <= 3834;
			WHEN "100101101011" => table_out <= 3834;
			WHEN "100101101100" => table_out <= 3834;
			WHEN "100101101101" => table_out <= 3834;
			WHEN "100101101110" => table_out <= 3834;
			WHEN "100101101111" => table_out <= 3835;
			WHEN "100101110000" => table_out <= 3835;
			WHEN "100101110001" => table_out <= 3835;
			WHEN "100101110010" => table_out <= 3835;
			WHEN "100101110011" => table_out <= 3835;
			WHEN "100101110100" => table_out <= 3836;
			WHEN "100101110101" => table_out <= 3836;
			WHEN "100101110110" => table_out <= 3836;
			WHEN "100101110111" => table_out <= 3836;
			WHEN "100101111000" => table_out <= 3836;
			WHEN "100101111001" => table_out <= 3837;
			WHEN "100101111010" => table_out <= 3837;
			WHEN "100101111011" => table_out <= 3837;
			WHEN "100101111100" => table_out <= 3837;
			WHEN "100101111101" => table_out <= 3837;
			WHEN "100101111110" => table_out <= 3838;
			WHEN "100101111111" => table_out <= 3838;
			WHEN "100110000000" => table_out <= 3838;
			WHEN "100110000001" => table_out <= 3838;
			WHEN "100110000010" => table_out <= 3838;
			WHEN "100110000011" => table_out <= 3839;
			WHEN "100110000100" => table_out <= 3839;
			WHEN "100110000101" => table_out <= 3839;
			WHEN "100110000110" => table_out <= 3839;
			WHEN "100110000111" => table_out <= 3839;
			WHEN "100110001000" => table_out <= 3840;
			WHEN "100110001001" => table_out <= 3840;
			WHEN "100110001010" => table_out <= 3840;
			WHEN "100110001011" => table_out <= 3840;
			WHEN "100110001100" => table_out <= 3840;
			WHEN "100110001101" => table_out <= 3841;
			WHEN "100110001110" => table_out <= 3841;
			WHEN "100110001111" => table_out <= 3841;
			WHEN "100110010000" => table_out <= 3841;
			WHEN "100110010001" => table_out <= 3841;
			WHEN "100110010010" => table_out <= 3842;
			WHEN "100110010011" => table_out <= 3842;
			WHEN "100110010100" => table_out <= 3842;
			WHEN "100110010101" => table_out <= 3842;
			WHEN "100110010110" => table_out <= 3842;
			WHEN "100110010111" => table_out <= 3843;
			WHEN "100110011000" => table_out <= 3843;
			WHEN "100110011001" => table_out <= 3843;
			WHEN "100110011010" => table_out <= 3843;
			WHEN "100110011011" => table_out <= 3843;
			WHEN "100110011100" => table_out <= 3844;
			WHEN "100110011101" => table_out <= 3844;
			WHEN "100110011110" => table_out <= 3844;
			WHEN "100110011111" => table_out <= 3844;
			WHEN "100110100000" => table_out <= 3844;
			WHEN "100110100001" => table_out <= 3845;
			WHEN "100110100010" => table_out <= 3845;
			WHEN "100110100011" => table_out <= 3845;
			WHEN "100110100100" => table_out <= 3845;
			WHEN "100110100101" => table_out <= 3845;
			WHEN "100110100110" => table_out <= 3846;
			WHEN "100110100111" => table_out <= 3846;
			WHEN "100110101000" => table_out <= 3846;
			WHEN "100110101001" => table_out <= 3846;
			WHEN "100110101010" => table_out <= 3846;
			WHEN "100110101011" => table_out <= 3847;
			WHEN "100110101100" => table_out <= 3847;
			WHEN "100110101101" => table_out <= 3847;
			WHEN "100110101110" => table_out <= 3847;
			WHEN "100110101111" => table_out <= 3847;
			WHEN "100110110000" => table_out <= 3848;
			WHEN "100110110001" => table_out <= 3848;
			WHEN "100110110010" => table_out <= 3848;
			WHEN "100110110011" => table_out <= 3848;
			WHEN "100110110100" => table_out <= 3848;
			WHEN "100110110101" => table_out <= 3849;
			WHEN "100110110110" => table_out <= 3849;
			WHEN "100110110111" => table_out <= 3849;
			WHEN "100110111000" => table_out <= 3849;
			WHEN "100110111001" => table_out <= 3849;
			WHEN "100110111010" => table_out <= 3850;
			WHEN "100110111011" => table_out <= 3850;
			WHEN "100110111100" => table_out <= 3850;
			WHEN "100110111101" => table_out <= 3850;
			WHEN "100110111110" => table_out <= 3850;
			WHEN "100110111111" => table_out <= 3851;
			WHEN "100111000000" => table_out <= 3851;
			WHEN "100111000001" => table_out <= 3851;
			WHEN "100111000010" => table_out <= 3851;
			WHEN "100111000011" => table_out <= 3851;
			WHEN "100111000100" => table_out <= 3852;
			WHEN "100111000101" => table_out <= 3852;
			WHEN "100111000110" => table_out <= 3852;
			WHEN "100111000111" => table_out <= 3852;
			WHEN "100111001000" => table_out <= 3852;
			WHEN "100111001001" => table_out <= 3853;
			WHEN "100111001010" => table_out <= 3853;
			WHEN "100111001011" => table_out <= 3853;
			WHEN "100111001100" => table_out <= 3853;
			WHEN "100111001101" => table_out <= 3853;
			WHEN "100111001110" => table_out <= 3854;
			WHEN "100111001111" => table_out <= 3854;
			WHEN "100111010000" => table_out <= 3854;
			WHEN "100111010001" => table_out <= 3854;
			WHEN "100111010010" => table_out <= 3854;
			WHEN "100111010011" => table_out <= 3855;
			WHEN "100111010100" => table_out <= 3855;
			WHEN "100111010101" => table_out <= 3855;
			WHEN "100111010110" => table_out <= 3855;
			WHEN "100111010111" => table_out <= 3855;
			WHEN "100111011000" => table_out <= 3856;
			WHEN "100111011001" => table_out <= 3856;
			WHEN "100111011010" => table_out <= 3856;
			WHEN "100111011011" => table_out <= 3856;
			WHEN "100111011100" => table_out <= 3856;
			WHEN "100111011101" => table_out <= 3857;
			WHEN "100111011110" => table_out <= 3857;
			WHEN "100111011111" => table_out <= 3857;
			WHEN "100111100000" => table_out <= 3857;
			WHEN "100111100001" => table_out <= 3857;
			WHEN "100111100010" => table_out <= 3857;
			WHEN "100111100011" => table_out <= 3858;
			WHEN "100111100100" => table_out <= 3858;
			WHEN "100111100101" => table_out <= 3858;
			WHEN "100111100110" => table_out <= 3858;
			WHEN "100111100111" => table_out <= 3858;
			WHEN "100111101000" => table_out <= 3859;
			WHEN "100111101001" => table_out <= 3859;
			WHEN "100111101010" => table_out <= 3859;
			WHEN "100111101011" => table_out <= 3859;
			WHEN "100111101100" => table_out <= 3859;
			WHEN "100111101101" => table_out <= 3860;
			WHEN "100111101110" => table_out <= 3860;
			WHEN "100111101111" => table_out <= 3860;
			WHEN "100111110000" => table_out <= 3860;
			WHEN "100111110001" => table_out <= 3860;
			WHEN "100111110010" => table_out <= 3861;
			WHEN "100111110011" => table_out <= 3861;
			WHEN "100111110100" => table_out <= 3861;
			WHEN "100111110101" => table_out <= 3861;
			WHEN "100111110110" => table_out <= 3861;
			WHEN "100111110111" => table_out <= 3862;
			WHEN "100111111000" => table_out <= 3862;
			WHEN "100111111001" => table_out <= 3862;
			WHEN "100111111010" => table_out <= 3862;
			WHEN "100111111011" => table_out <= 3862;
			WHEN "100111111100" => table_out <= 3863;
			WHEN "100111111101" => table_out <= 3863;
			WHEN "100111111110" => table_out <= 3863;
			WHEN "100111111111" => table_out <= 3863;
			WHEN "101000000000" => table_out <= 3863;
			WHEN "101000000001" => table_out <= 3863;
			WHEN "101000000010" => table_out <= 3864;
			WHEN "101000000011" => table_out <= 3864;
			WHEN "101000000100" => table_out <= 3864;
			WHEN "101000000101" => table_out <= 3864;
			WHEN "101000000110" => table_out <= 3864;
			WHEN "101000000111" => table_out <= 3865;
			WHEN "101000001000" => table_out <= 3865;
			WHEN "101000001001" => table_out <= 3865;
			WHEN "101000001010" => table_out <= 3865;
			WHEN "101000001011" => table_out <= 3865;
			WHEN "101000001100" => table_out <= 3866;
			WHEN "101000001101" => table_out <= 3866;
			WHEN "101000001110" => table_out <= 3866;
			WHEN "101000001111" => table_out <= 3866;
			WHEN "101000010000" => table_out <= 3866;
			WHEN "101000010001" => table_out <= 3867;
			WHEN "101000010010" => table_out <= 3867;
			WHEN "101000010011" => table_out <= 3867;
			WHEN "101000010100" => table_out <= 3867;
			WHEN "101000010101" => table_out <= 3867;
			WHEN "101000010110" => table_out <= 3867;
			WHEN "101000010111" => table_out <= 3868;
			WHEN "101000011000" => table_out <= 3868;
			WHEN "101000011001" => table_out <= 3868;
			WHEN "101000011010" => table_out <= 3868;
			WHEN "101000011011" => table_out <= 3868;
			WHEN "101000011100" => table_out <= 3869;
			WHEN "101000011101" => table_out <= 3869;
			WHEN "101000011110" => table_out <= 3869;
			WHEN "101000011111" => table_out <= 3869;
			WHEN "101000100000" => table_out <= 3869;
			WHEN "101000100001" => table_out <= 3870;
			WHEN "101000100010" => table_out <= 3870;
			WHEN "101000100011" => table_out <= 3870;
			WHEN "101000100100" => table_out <= 3870;
			WHEN "101000100101" => table_out <= 3870;
			WHEN "101000100110" => table_out <= 3871;
			WHEN "101000100111" => table_out <= 3871;
			WHEN "101000101000" => table_out <= 3871;
			WHEN "101000101001" => table_out <= 3871;
			WHEN "101000101010" => table_out <= 3871;
			WHEN "101000101011" => table_out <= 3871;
			WHEN "101000101100" => table_out <= 3872;
			WHEN "101000101101" => table_out <= 3872;
			WHEN "101000101110" => table_out <= 3872;
			WHEN "101000101111" => table_out <= 3872;
			WHEN "101000110000" => table_out <= 3872;
			WHEN "101000110001" => table_out <= 3873;
			WHEN "101000110010" => table_out <= 3873;
			WHEN "101000110011" => table_out <= 3873;
			WHEN "101000110100" => table_out <= 3873;
			WHEN "101000110101" => table_out <= 3873;
			WHEN "101000110110" => table_out <= 3874;
			WHEN "101000110111" => table_out <= 3874;
			WHEN "101000111000" => table_out <= 3874;
			WHEN "101000111001" => table_out <= 3874;
			WHEN "101000111010" => table_out <= 3874;
			WHEN "101000111011" => table_out <= 3874;
			WHEN "101000111100" => table_out <= 3875;
			WHEN "101000111101" => table_out <= 3875;
			WHEN "101000111110" => table_out <= 3875;
			WHEN "101000111111" => table_out <= 3875;
			WHEN "101001000000" => table_out <= 3875;
			WHEN "101001000001" => table_out <= 3876;
			WHEN "101001000010" => table_out <= 3876;
			WHEN "101001000011" => table_out <= 3876;
			WHEN "101001000100" => table_out <= 3876;
			WHEN "101001000101" => table_out <= 3876;
			WHEN "101001000110" => table_out <= 3877;
			WHEN "101001000111" => table_out <= 3877;
			WHEN "101001001000" => table_out <= 3877;
			WHEN "101001001001" => table_out <= 3877;
			WHEN "101001001010" => table_out <= 3877;
			WHEN "101001001011" => table_out <= 3877;
			WHEN "101001001100" => table_out <= 3878;
			WHEN "101001001101" => table_out <= 3878;
			WHEN "101001001110" => table_out <= 3878;
			WHEN "101001001111" => table_out <= 3878;
			WHEN "101001010000" => table_out <= 3878;
			WHEN "101001010001" => table_out <= 3879;
			WHEN "101001010010" => table_out <= 3879;
			WHEN "101001010011" => table_out <= 3879;
			WHEN "101001010100" => table_out <= 3879;
			WHEN "101001010101" => table_out <= 3879;
			WHEN "101001010110" => table_out <= 3880;
			WHEN "101001010111" => table_out <= 3880;
			WHEN "101001011000" => table_out <= 3880;
			WHEN "101001011001" => table_out <= 3880;
			WHEN "101001011010" => table_out <= 3880;
			WHEN "101001011011" => table_out <= 3880;
			WHEN "101001011100" => table_out <= 3881;
			WHEN "101001011101" => table_out <= 3881;
			WHEN "101001011110" => table_out <= 3881;
			WHEN "101001011111" => table_out <= 3881;
			WHEN "101001100000" => table_out <= 3881;
			WHEN "101001100001" => table_out <= 3882;
			WHEN "101001100010" => table_out <= 3882;
			WHEN "101001100011" => table_out <= 3882;
			WHEN "101001100100" => table_out <= 3882;
			WHEN "101001100101" => table_out <= 3882;
			WHEN "101001100110" => table_out <= 3883;
			WHEN "101001100111" => table_out <= 3883;
			WHEN "101001101000" => table_out <= 3883;
			WHEN "101001101001" => table_out <= 3883;
			WHEN "101001101010" => table_out <= 3883;
			WHEN "101001101011" => table_out <= 3883;
			WHEN "101001101100" => table_out <= 3884;
			WHEN "101001101101" => table_out <= 3884;
			WHEN "101001101110" => table_out <= 3884;
			WHEN "101001101111" => table_out <= 3884;
			WHEN "101001110000" => table_out <= 3884;
			WHEN "101001110001" => table_out <= 3885;
			WHEN "101001110010" => table_out <= 3885;
			WHEN "101001110011" => table_out <= 3885;
			WHEN "101001110100" => table_out <= 3885;
			WHEN "101001110101" => table_out <= 3885;
			WHEN "101001110110" => table_out <= 3885;
			WHEN "101001110111" => table_out <= 3886;
			WHEN "101001111000" => table_out <= 3886;
			WHEN "101001111001" => table_out <= 3886;
			WHEN "101001111010" => table_out <= 3886;
			WHEN "101001111011" => table_out <= 3886;
			WHEN "101001111100" => table_out <= 3887;
			WHEN "101001111101" => table_out <= 3887;
			WHEN "101001111110" => table_out <= 3887;
			WHEN "101001111111" => table_out <= 3887;
			WHEN "101010000000" => table_out <= 3887;
			WHEN "101010000001" => table_out <= 3887;
			WHEN "101010000010" => table_out <= 3888;
			WHEN "101010000011" => table_out <= 3888;
			WHEN "101010000100" => table_out <= 3888;
			WHEN "101010000101" => table_out <= 3888;
			WHEN "101010000110" => table_out <= 3888;
			WHEN "101010000111" => table_out <= 3889;
			WHEN "101010001000" => table_out <= 3889;
			WHEN "101010001001" => table_out <= 3889;
			WHEN "101010001010" => table_out <= 3889;
			WHEN "101010001011" => table_out <= 3889;
			WHEN "101010001100" => table_out <= 3889;
			WHEN "101010001101" => table_out <= 3890;
			WHEN "101010001110" => table_out <= 3890;
			WHEN "101010001111" => table_out <= 3890;
			WHEN "101010010000" => table_out <= 3890;
			WHEN "101010010001" => table_out <= 3890;
			WHEN "101010010010" => table_out <= 3891;
			WHEN "101010010011" => table_out <= 3891;
			WHEN "101010010100" => table_out <= 3891;
			WHEN "101010010101" => table_out <= 3891;
			WHEN "101010010110" => table_out <= 3891;
			WHEN "101010010111" => table_out <= 3891;
			WHEN "101010011000" => table_out <= 3892;
			WHEN "101010011001" => table_out <= 3892;
			WHEN "101010011010" => table_out <= 3892;
			WHEN "101010011011" => table_out <= 3892;
			WHEN "101010011100" => table_out <= 3892;
			WHEN "101010011101" => table_out <= 3893;
			WHEN "101010011110" => table_out <= 3893;
			WHEN "101010011111" => table_out <= 3893;
			WHEN "101010100000" => table_out <= 3893;
			WHEN "101010100001" => table_out <= 3893;
			WHEN "101010100010" => table_out <= 3893;
			WHEN "101010100011" => table_out <= 3894;
			WHEN "101010100100" => table_out <= 3894;
			WHEN "101010100101" => table_out <= 3894;
			WHEN "101010100110" => table_out <= 3894;
			WHEN "101010100111" => table_out <= 3894;
			WHEN "101010101000" => table_out <= 3895;
			WHEN "101010101001" => table_out <= 3895;
			WHEN "101010101010" => table_out <= 3895;
			WHEN "101010101011" => table_out <= 3895;
			WHEN "101010101100" => table_out <= 3895;
			WHEN "101010101101" => table_out <= 3895;
			WHEN "101010101110" => table_out <= 3896;
			WHEN "101010101111" => table_out <= 3896;
			WHEN "101010110000" => table_out <= 3896;
			WHEN "101010110001" => table_out <= 3896;
			WHEN "101010110010" => table_out <= 3896;
			WHEN "101010110011" => table_out <= 3897;
			WHEN "101010110100" => table_out <= 3897;
			WHEN "101010110101" => table_out <= 3897;
			WHEN "101010110110" => table_out <= 3897;
			WHEN "101010110111" => table_out <= 3897;
			WHEN "101010111000" => table_out <= 3897;
			WHEN "101010111001" => table_out <= 3898;
			WHEN "101010111010" => table_out <= 3898;
			WHEN "101010111011" => table_out <= 3898;
			WHEN "101010111100" => table_out <= 3898;
			WHEN "101010111101" => table_out <= 3898;
			WHEN "101010111110" => table_out <= 3899;
			WHEN "101010111111" => table_out <= 3899;
			WHEN "101011000000" => table_out <= 3899;
			WHEN "101011000001" => table_out <= 3899;
			WHEN "101011000010" => table_out <= 3899;
			WHEN "101011000011" => table_out <= 3899;
			WHEN "101011000100" => table_out <= 3900;
			WHEN "101011000101" => table_out <= 3900;
			WHEN "101011000110" => table_out <= 3900;
			WHEN "101011000111" => table_out <= 3900;
			WHEN "101011001000" => table_out <= 3900;
			WHEN "101011001001" => table_out <= 3900;
			WHEN "101011001010" => table_out <= 3901;
			WHEN "101011001011" => table_out <= 3901;
			WHEN "101011001100" => table_out <= 3901;
			WHEN "101011001101" => table_out <= 3901;
			WHEN "101011001110" => table_out <= 3901;
			WHEN "101011001111" => table_out <= 3902;
			WHEN "101011010000" => table_out <= 3902;
			WHEN "101011010001" => table_out <= 3902;
			WHEN "101011010010" => table_out <= 3902;
			WHEN "101011010011" => table_out <= 3902;
			WHEN "101011010100" => table_out <= 3902;
			WHEN "101011010101" => table_out <= 3903;
			WHEN "101011010110" => table_out <= 3903;
			WHEN "101011010111" => table_out <= 3903;
			WHEN "101011011000" => table_out <= 3903;
			WHEN "101011011001" => table_out <= 3903;
			WHEN "101011011010" => table_out <= 3904;
			WHEN "101011011011" => table_out <= 3904;
			WHEN "101011011100" => table_out <= 3904;
			WHEN "101011011101" => table_out <= 3904;
			WHEN "101011011110" => table_out <= 3904;
			WHEN "101011011111" => table_out <= 3904;
			WHEN "101011100000" => table_out <= 3905;
			WHEN "101011100001" => table_out <= 3905;
			WHEN "101011100010" => table_out <= 3905;
			WHEN "101011100011" => table_out <= 3905;
			WHEN "101011100100" => table_out <= 3905;
			WHEN "101011100101" => table_out <= 3905;
			WHEN "101011100110" => table_out <= 3906;
			WHEN "101011100111" => table_out <= 3906;
			WHEN "101011101000" => table_out <= 3906;
			WHEN "101011101001" => table_out <= 3906;
			WHEN "101011101010" => table_out <= 3906;
			WHEN "101011101011" => table_out <= 3907;
			WHEN "101011101100" => table_out <= 3907;
			WHEN "101011101101" => table_out <= 3907;
			WHEN "101011101110" => table_out <= 3907;
			WHEN "101011101111" => table_out <= 3907;
			WHEN "101011110000" => table_out <= 3907;
			WHEN "101011110001" => table_out <= 3908;
			WHEN "101011110010" => table_out <= 3908;
			WHEN "101011110011" => table_out <= 3908;
			WHEN "101011110100" => table_out <= 3908;
			WHEN "101011110101" => table_out <= 3908;
			WHEN "101011110110" => table_out <= 3908;
			WHEN "101011110111" => table_out <= 3909;
			WHEN "101011111000" => table_out <= 3909;
			WHEN "101011111001" => table_out <= 3909;
			WHEN "101011111010" => table_out <= 3909;
			WHEN "101011111011" => table_out <= 3909;
			WHEN "101011111100" => table_out <= 3909;
			WHEN "101011111101" => table_out <= 3910;
			WHEN "101011111110" => table_out <= 3910;
			WHEN "101011111111" => table_out <= 3910;
			WHEN "101100000000" => table_out <= 3910;
			WHEN "101100000001" => table_out <= 3910;
			WHEN "101100000010" => table_out <= 3911;
			WHEN "101100000011" => table_out <= 3911;
			WHEN "101100000100" => table_out <= 3911;
			WHEN "101100000101" => table_out <= 3911;
			WHEN "101100000110" => table_out <= 3911;
			WHEN "101100000111" => table_out <= 3911;
			WHEN "101100001000" => table_out <= 3912;
			WHEN "101100001001" => table_out <= 3912;
			WHEN "101100001010" => table_out <= 3912;
			WHEN "101100001011" => table_out <= 3912;
			WHEN "101100001100" => table_out <= 3912;
			WHEN "101100001101" => table_out <= 3912;
			WHEN "101100001110" => table_out <= 3913;
			WHEN "101100001111" => table_out <= 3913;
			WHEN "101100010000" => table_out <= 3913;
			WHEN "101100010001" => table_out <= 3913;
			WHEN "101100010010" => table_out <= 3913;
			WHEN "101100010011" => table_out <= 3914;
			WHEN "101100010100" => table_out <= 3914;
			WHEN "101100010101" => table_out <= 3914;
			WHEN "101100010110" => table_out <= 3914;
			WHEN "101100010111" => table_out <= 3914;
			WHEN "101100011000" => table_out <= 3914;
			WHEN "101100011001" => table_out <= 3915;
			WHEN "101100011010" => table_out <= 3915;
			WHEN "101100011011" => table_out <= 3915;
			WHEN "101100011100" => table_out <= 3915;
			WHEN "101100011101" => table_out <= 3915;
			WHEN "101100011110" => table_out <= 3915;
			WHEN "101100011111" => table_out <= 3916;
			WHEN "101100100000" => table_out <= 3916;
			WHEN "101100100001" => table_out <= 3916;
			WHEN "101100100010" => table_out <= 3916;
			WHEN "101100100011" => table_out <= 3916;
			WHEN "101100100100" => table_out <= 3916;
			WHEN "101100100101" => table_out <= 3917;
			WHEN "101100100110" => table_out <= 3917;
			WHEN "101100100111" => table_out <= 3917;
			WHEN "101100101000" => table_out <= 3917;
			WHEN "101100101001" => table_out <= 3917;
			WHEN "101100101010" => table_out <= 3917;
			WHEN "101100101011" => table_out <= 3918;
			WHEN "101100101100" => table_out <= 3918;
			WHEN "101100101101" => table_out <= 3918;
			WHEN "101100101110" => table_out <= 3918;
			WHEN "101100101111" => table_out <= 3918;
			WHEN "101100110000" => table_out <= 3919;
			WHEN "101100110001" => table_out <= 3919;
			WHEN "101100110010" => table_out <= 3919;
			WHEN "101100110011" => table_out <= 3919;
			WHEN "101100110100" => table_out <= 3919;
			WHEN "101100110101" => table_out <= 3919;
			WHEN "101100110110" => table_out <= 3920;
			WHEN "101100110111" => table_out <= 3920;
			WHEN "101100111000" => table_out <= 3920;
			WHEN "101100111001" => table_out <= 3920;
			WHEN "101100111010" => table_out <= 3920;
			WHEN "101100111011" => table_out <= 3920;
			WHEN "101100111100" => table_out <= 3921;
			WHEN "101100111101" => table_out <= 3921;
			WHEN "101100111110" => table_out <= 3921;
			WHEN "101100111111" => table_out <= 3921;
			WHEN "101101000000" => table_out <= 3921;
			WHEN "101101000001" => table_out <= 3921;
			WHEN "101101000010" => table_out <= 3922;
			WHEN "101101000011" => table_out <= 3922;
			WHEN "101101000100" => table_out <= 3922;
			WHEN "101101000101" => table_out <= 3922;
			WHEN "101101000110" => table_out <= 3922;
			WHEN "101101000111" => table_out <= 3922;
			WHEN "101101001000" => table_out <= 3923;
			WHEN "101101001001" => table_out <= 3923;
			WHEN "101101001010" => table_out <= 3923;
			WHEN "101101001011" => table_out <= 3923;
			WHEN "101101001100" => table_out <= 3923;
			WHEN "101101001101" => table_out <= 3923;
			WHEN "101101001110" => table_out <= 3924;
			WHEN "101101001111" => table_out <= 3924;
			WHEN "101101010000" => table_out <= 3924;
			WHEN "101101010001" => table_out <= 3924;
			WHEN "101101010010" => table_out <= 3924;
			WHEN "101101010011" => table_out <= 3924;
			WHEN "101101010100" => table_out <= 3925;
			WHEN "101101010101" => table_out <= 3925;
			WHEN "101101010110" => table_out <= 3925;
			WHEN "101101010111" => table_out <= 3925;
			WHEN "101101011000" => table_out <= 3925;
			WHEN "101101011001" => table_out <= 3926;
			WHEN "101101011010" => table_out <= 3926;
			WHEN "101101011011" => table_out <= 3926;
			WHEN "101101011100" => table_out <= 3926;
			WHEN "101101011101" => table_out <= 3926;
			WHEN "101101011110" => table_out <= 3926;
			WHEN "101101011111" => table_out <= 3927;
			WHEN "101101100000" => table_out <= 3927;
			WHEN "101101100001" => table_out <= 3927;
			WHEN "101101100010" => table_out <= 3927;
			WHEN "101101100011" => table_out <= 3927;
			WHEN "101101100100" => table_out <= 3927;
			WHEN "101101100101" => table_out <= 3928;
			WHEN "101101100110" => table_out <= 3928;
			WHEN "101101100111" => table_out <= 3928;
			WHEN "101101101000" => table_out <= 3928;
			WHEN "101101101001" => table_out <= 3928;
			WHEN "101101101010" => table_out <= 3928;
			WHEN "101101101011" => table_out <= 3929;
			WHEN "101101101100" => table_out <= 3929;
			WHEN "101101101101" => table_out <= 3929;
			WHEN "101101101110" => table_out <= 3929;
			WHEN "101101101111" => table_out <= 3929;
			WHEN "101101110000" => table_out <= 3929;
			WHEN "101101110001" => table_out <= 3930;
			WHEN "101101110010" => table_out <= 3930;
			WHEN "101101110011" => table_out <= 3930;
			WHEN "101101110100" => table_out <= 3930;
			WHEN "101101110101" => table_out <= 3930;
			WHEN "101101110110" => table_out <= 3930;
			WHEN "101101110111" => table_out <= 3931;
			WHEN "101101111000" => table_out <= 3931;
			WHEN "101101111001" => table_out <= 3931;
			WHEN "101101111010" => table_out <= 3931;
			WHEN "101101111011" => table_out <= 3931;
			WHEN "101101111100" => table_out <= 3931;
			WHEN "101101111101" => table_out <= 3932;
			WHEN "101101111110" => table_out <= 3932;
			WHEN "101101111111" => table_out <= 3932;
			WHEN "101110000000" => table_out <= 3932;
			WHEN "101110000001" => table_out <= 3932;
			WHEN "101110000010" => table_out <= 3932;
			WHEN "101110000011" => table_out <= 3933;
			WHEN "101110000100" => table_out <= 3933;
			WHEN "101110000101" => table_out <= 3933;
			WHEN "101110000110" => table_out <= 3933;
			WHEN "101110000111" => table_out <= 3933;
			WHEN "101110001000" => table_out <= 3933;
			WHEN "101110001001" => table_out <= 3934;
			WHEN "101110001010" => table_out <= 3934;
			WHEN "101110001011" => table_out <= 3934;
			WHEN "101110001100" => table_out <= 3934;
			WHEN "101110001101" => table_out <= 3934;
			WHEN "101110001110" => table_out <= 3934;
			WHEN "101110001111" => table_out <= 3935;
			WHEN "101110010000" => table_out <= 3935;
			WHEN "101110010001" => table_out <= 3935;
			WHEN "101110010010" => table_out <= 3935;
			WHEN "101110010011" => table_out <= 3935;
			WHEN "101110010100" => table_out <= 3935;
			WHEN "101110010101" => table_out <= 3936;
			WHEN "101110010110" => table_out <= 3936;
			WHEN "101110010111" => table_out <= 3936;
			WHEN "101110011000" => table_out <= 3936;
			WHEN "101110011001" => table_out <= 3936;
			WHEN "101110011010" => table_out <= 3936;
			WHEN "101110011011" => table_out <= 3937;
			WHEN "101110011100" => table_out <= 3937;
			WHEN "101110011101" => table_out <= 3937;
			WHEN "101110011110" => table_out <= 3937;
			WHEN "101110011111" => table_out <= 3937;
			WHEN "101110100000" => table_out <= 3937;
			WHEN "101110100001" => table_out <= 3938;
			WHEN "101110100010" => table_out <= 3938;
			WHEN "101110100011" => table_out <= 3938;
			WHEN "101110100100" => table_out <= 3938;
			WHEN "101110100101" => table_out <= 3938;
			WHEN "101110100110" => table_out <= 3938;
			WHEN "101110100111" => table_out <= 3939;
			WHEN "101110101000" => table_out <= 3939;
			WHEN "101110101001" => table_out <= 3939;
			WHEN "101110101010" => table_out <= 3939;
			WHEN "101110101011" => table_out <= 3939;
			WHEN "101110101100" => table_out <= 3939;
			WHEN "101110101101" => table_out <= 3940;
			WHEN "101110101110" => table_out <= 3940;
			WHEN "101110101111" => table_out <= 3940;
			WHEN "101110110000" => table_out <= 3940;
			WHEN "101110110001" => table_out <= 3940;
			WHEN "101110110010" => table_out <= 3940;
			WHEN "101110110011" => table_out <= 3941;
			WHEN "101110110100" => table_out <= 3941;
			WHEN "101110110101" => table_out <= 3941;
			WHEN "101110110110" => table_out <= 3941;
			WHEN "101110110111" => table_out <= 3941;
			WHEN "101110111000" => table_out <= 3941;
			WHEN "101110111001" => table_out <= 3942;
			WHEN "101110111010" => table_out <= 3942;
			WHEN "101110111011" => table_out <= 3942;
			WHEN "101110111100" => table_out <= 3942;
			WHEN "101110111101" => table_out <= 3942;
			WHEN "101110111110" => table_out <= 3942;
			WHEN "101110111111" => table_out <= 3942;
			WHEN "101111000000" => table_out <= 3943;
			WHEN "101111000001" => table_out <= 3943;
			WHEN "101111000010" => table_out <= 3943;
			WHEN "101111000011" => table_out <= 3943;
			WHEN "101111000100" => table_out <= 3943;
			WHEN "101111000101" => table_out <= 3943;
			WHEN "101111000110" => table_out <= 3944;
			WHEN "101111000111" => table_out <= 3944;
			WHEN "101111001000" => table_out <= 3944;
			WHEN "101111001001" => table_out <= 3944;
			WHEN "101111001010" => table_out <= 3944;
			WHEN "101111001011" => table_out <= 3944;
			WHEN "101111001100" => table_out <= 3945;
			WHEN "101111001101" => table_out <= 3945;
			WHEN "101111001110" => table_out <= 3945;
			WHEN "101111001111" => table_out <= 3945;
			WHEN "101111010000" => table_out <= 3945;
			WHEN "101111010001" => table_out <= 3945;
			WHEN "101111010010" => table_out <= 3946;
			WHEN "101111010011" => table_out <= 3946;
			WHEN "101111010100" => table_out <= 3946;
			WHEN "101111010101" => table_out <= 3946;
			WHEN "101111010110" => table_out <= 3946;
			WHEN "101111010111" => table_out <= 3946;
			WHEN "101111011000" => table_out <= 3947;
			WHEN "101111011001" => table_out <= 3947;
			WHEN "101111011010" => table_out <= 3947;
			WHEN "101111011011" => table_out <= 3947;
			WHEN "101111011100" => table_out <= 3947;
			WHEN "101111011101" => table_out <= 3947;
			WHEN "101111011110" => table_out <= 3948;
			WHEN "101111011111" => table_out <= 3948;
			WHEN "101111100000" => table_out <= 3948;
			WHEN "101111100001" => table_out <= 3948;
			WHEN "101111100010" => table_out <= 3948;
			WHEN "101111100011" => table_out <= 3948;
			WHEN "101111100100" => table_out <= 3949;
			WHEN "101111100101" => table_out <= 3949;
			WHEN "101111100110" => table_out <= 3949;
			WHEN "101111100111" => table_out <= 3949;
			WHEN "101111101000" => table_out <= 3949;
			WHEN "101111101001" => table_out <= 3949;
			WHEN "101111101010" => table_out <= 3949;
			WHEN "101111101011" => table_out <= 3950;
			WHEN "101111101100" => table_out <= 3950;
			WHEN "101111101101" => table_out <= 3950;
			WHEN "101111101110" => table_out <= 3950;
			WHEN "101111101111" => table_out <= 3950;
			WHEN "101111110000" => table_out <= 3950;
			WHEN "101111110001" => table_out <= 3951;
			WHEN "101111110010" => table_out <= 3951;
			WHEN "101111110011" => table_out <= 3951;
			WHEN "101111110100" => table_out <= 3951;
			WHEN "101111110101" => table_out <= 3951;
			WHEN "101111110110" => table_out <= 3951;
			WHEN "101111110111" => table_out <= 3952;
			WHEN "101111111000" => table_out <= 3952;
			WHEN "101111111001" => table_out <= 3952;
			WHEN "101111111010" => table_out <= 3952;
			WHEN "101111111011" => table_out <= 3952;
			WHEN "101111111100" => table_out <= 3952;
			WHEN "101111111101" => table_out <= 3953;
			WHEN "101111111110" => table_out <= 3953;
			WHEN "101111111111" => table_out <= 3953;
			WHEN "110000000000" => table_out <= 3953;
			WHEN "110000000001" => table_out <= 3953;
			WHEN "110000000010" => table_out <= 3953;
			WHEN "110000000011" => table_out <= 3953;
			WHEN "110000000100" => table_out <= 3954;
			WHEN "110000000101" => table_out <= 3954;
			WHEN "110000000110" => table_out <= 3954;
			WHEN "110000000111" => table_out <= 3954;
			WHEN "110000001000" => table_out <= 3954;
			WHEN "110000001001" => table_out <= 3954;
			WHEN "110000001010" => table_out <= 3955;
			WHEN "110000001011" => table_out <= 3955;
			WHEN "110000001100" => table_out <= 3955;
			WHEN "110000001101" => table_out <= 3955;
			WHEN "110000001110" => table_out <= 3955;
			WHEN "110000001111" => table_out <= 3955;
			WHEN "110000010000" => table_out <= 3956;
			WHEN "110000010001" => table_out <= 3956;
			WHEN "110000010010" => table_out <= 3956;
			WHEN "110000010011" => table_out <= 3956;
			WHEN "110000010100" => table_out <= 3956;
			WHEN "110000010101" => table_out <= 3956;
			WHEN "110000010110" => table_out <= 3957;
			WHEN "110000010111" => table_out <= 3957;
			WHEN "110000011000" => table_out <= 3957;
			WHEN "110000011001" => table_out <= 3957;
			WHEN "110000011010" => table_out <= 3957;
			WHEN "110000011011" => table_out <= 3957;
			WHEN "110000011100" => table_out <= 3957;
			WHEN "110000011101" => table_out <= 3958;
			WHEN "110000011110" => table_out <= 3958;
			WHEN "110000011111" => table_out <= 3958;
			WHEN "110000100000" => table_out <= 3958;
			WHEN "110000100001" => table_out <= 3958;
			WHEN "110000100010" => table_out <= 3958;
			WHEN "110000100011" => table_out <= 3959;
			WHEN "110000100100" => table_out <= 3959;
			WHEN "110000100101" => table_out <= 3959;
			WHEN "110000100110" => table_out <= 3959;
			WHEN "110000100111" => table_out <= 3959;
			WHEN "110000101000" => table_out <= 3959;
			WHEN "110000101001" => table_out <= 3960;
			WHEN "110000101010" => table_out <= 3960;
			WHEN "110000101011" => table_out <= 3960;
			WHEN "110000101100" => table_out <= 3960;
			WHEN "110000101101" => table_out <= 3960;
			WHEN "110000101110" => table_out <= 3960;
			WHEN "110000101111" => table_out <= 3960;
			WHEN "110000110000" => table_out <= 3961;
			WHEN "110000110001" => table_out <= 3961;
			WHEN "110000110010" => table_out <= 3961;
			WHEN "110000110011" => table_out <= 3961;
			WHEN "110000110100" => table_out <= 3961;
			WHEN "110000110101" => table_out <= 3961;
			WHEN "110000110110" => table_out <= 3962;
			WHEN "110000110111" => table_out <= 3962;
			WHEN "110000111000" => table_out <= 3962;
			WHEN "110000111001" => table_out <= 3962;
			WHEN "110000111010" => table_out <= 3962;
			WHEN "110000111011" => table_out <= 3962;
			WHEN "110000111100" => table_out <= 3963;
			WHEN "110000111101" => table_out <= 3963;
			WHEN "110000111110" => table_out <= 3963;
			WHEN "110000111111" => table_out <= 3963;
			WHEN "110001000000" => table_out <= 3963;
			WHEN "110001000001" => table_out <= 3963;
			WHEN "110001000010" => table_out <= 3963;
			WHEN "110001000011" => table_out <= 3964;
			WHEN "110001000100" => table_out <= 3964;
			WHEN "110001000101" => table_out <= 3964;
			WHEN "110001000110" => table_out <= 3964;
			WHEN "110001000111" => table_out <= 3964;
			WHEN "110001001000" => table_out <= 3964;
			WHEN "110001001001" => table_out <= 3965;
			WHEN "110001001010" => table_out <= 3965;
			WHEN "110001001011" => table_out <= 3965;
			WHEN "110001001100" => table_out <= 3965;
			WHEN "110001001101" => table_out <= 3965;
			WHEN "110001001110" => table_out <= 3965;
			WHEN "110001001111" => table_out <= 3966;
			WHEN "110001010000" => table_out <= 3966;
			WHEN "110001010001" => table_out <= 3966;
			WHEN "110001010010" => table_out <= 3966;
			WHEN "110001010011" => table_out <= 3966;
			WHEN "110001010100" => table_out <= 3966;
			WHEN "110001010101" => table_out <= 3966;
			WHEN "110001010110" => table_out <= 3967;
			WHEN "110001010111" => table_out <= 3967;
			WHEN "110001011000" => table_out <= 3967;
			WHEN "110001011001" => table_out <= 3967;
			WHEN "110001011010" => table_out <= 3967;
			WHEN "110001011011" => table_out <= 3967;
			WHEN "110001011100" => table_out <= 3968;
			WHEN "110001011101" => table_out <= 3968;
			WHEN "110001011110" => table_out <= 3968;
			WHEN "110001011111" => table_out <= 3968;
			WHEN "110001100000" => table_out <= 3968;
			WHEN "110001100001" => table_out <= 3968;
			WHEN "110001100010" => table_out <= 3968;
			WHEN "110001100011" => table_out <= 3969;
			WHEN "110001100100" => table_out <= 3969;
			WHEN "110001100101" => table_out <= 3969;
			WHEN "110001100110" => table_out <= 3969;
			WHEN "110001100111" => table_out <= 3969;
			WHEN "110001101000" => table_out <= 3969;
			WHEN "110001101001" => table_out <= 3970;
			WHEN "110001101010" => table_out <= 3970;
			WHEN "110001101011" => table_out <= 3970;
			WHEN "110001101100" => table_out <= 3970;
			WHEN "110001101101" => table_out <= 3970;
			WHEN "110001101110" => table_out <= 3970;
			WHEN "110001101111" => table_out <= 3970;
			WHEN "110001110000" => table_out <= 3971;
			WHEN "110001110001" => table_out <= 3971;
			WHEN "110001110010" => table_out <= 3971;
			WHEN "110001110011" => table_out <= 3971;
			WHEN "110001110100" => table_out <= 3971;
			WHEN "110001110101" => table_out <= 3971;
			WHEN "110001110110" => table_out <= 3972;
			WHEN "110001110111" => table_out <= 3972;
			WHEN "110001111000" => table_out <= 3972;
			WHEN "110001111001" => table_out <= 3972;
			WHEN "110001111010" => table_out <= 3972;
			WHEN "110001111011" => table_out <= 3972;
			WHEN "110001111100" => table_out <= 3972;
			WHEN "110001111101" => table_out <= 3973;
			WHEN "110001111110" => table_out <= 3973;
			WHEN "110001111111" => table_out <= 3973;
			WHEN "110010000000" => table_out <= 3973;
			WHEN "110010000001" => table_out <= 3973;
			WHEN "110010000010" => table_out <= 3973;
			WHEN "110010000011" => table_out <= 3974;
			WHEN "110010000100" => table_out <= 3974;
			WHEN "110010000101" => table_out <= 3974;
			WHEN "110010000110" => table_out <= 3974;
			WHEN "110010000111" => table_out <= 3974;
			WHEN "110010001000" => table_out <= 3974;
			WHEN "110010001001" => table_out <= 3974;
			WHEN "110010001010" => table_out <= 3975;
			WHEN "110010001011" => table_out <= 3975;
			WHEN "110010001100" => table_out <= 3975;
			WHEN "110010001101" => table_out <= 3975;
			WHEN "110010001110" => table_out <= 3975;
			WHEN "110010001111" => table_out <= 3975;
			WHEN "110010010000" => table_out <= 3976;
			WHEN "110010010001" => table_out <= 3976;
			WHEN "110010010010" => table_out <= 3976;
			WHEN "110010010011" => table_out <= 3976;
			WHEN "110010010100" => table_out <= 3976;
			WHEN "110010010101" => table_out <= 3976;
			WHEN "110010010110" => table_out <= 3976;
			WHEN "110010010111" => table_out <= 3977;
			WHEN "110010011000" => table_out <= 3977;
			WHEN "110010011001" => table_out <= 3977;
			WHEN "110010011010" => table_out <= 3977;
			WHEN "110010011011" => table_out <= 3977;
			WHEN "110010011100" => table_out <= 3977;
			WHEN "110010011101" => table_out <= 3978;
			WHEN "110010011110" => table_out <= 3978;
			WHEN "110010011111" => table_out <= 3978;
			WHEN "110010100000" => table_out <= 3978;
			WHEN "110010100001" => table_out <= 3978;
			WHEN "110010100010" => table_out <= 3978;
			WHEN "110010100011" => table_out <= 3978;
			WHEN "110010100100" => table_out <= 3979;
			WHEN "110010100101" => table_out <= 3979;
			WHEN "110010100110" => table_out <= 3979;
			WHEN "110010100111" => table_out <= 3979;
			WHEN "110010101000" => table_out <= 3979;
			WHEN "110010101001" => table_out <= 3979;
			WHEN "110010101010" => table_out <= 3980;
			WHEN "110010101011" => table_out <= 3980;
			WHEN "110010101100" => table_out <= 3980;
			WHEN "110010101101" => table_out <= 3980;
			WHEN "110010101110" => table_out <= 3980;
			WHEN "110010101111" => table_out <= 3980;
			WHEN "110010110000" => table_out <= 3980;
			WHEN "110010110001" => table_out <= 3981;
			WHEN "110010110010" => table_out <= 3981;
			WHEN "110010110011" => table_out <= 3981;
			WHEN "110010110100" => table_out <= 3981;
			WHEN "110010110101" => table_out <= 3981;
			WHEN "110010110110" => table_out <= 3981;
			WHEN "110010110111" => table_out <= 3982;
			WHEN "110010111000" => table_out <= 3982;
			WHEN "110010111001" => table_out <= 3982;
			WHEN "110010111010" => table_out <= 3982;
			WHEN "110010111011" => table_out <= 3982;
			WHEN "110010111100" => table_out <= 3982;
			WHEN "110010111101" => table_out <= 3982;
			WHEN "110010111110" => table_out <= 3983;
			WHEN "110010111111" => table_out <= 3983;
			WHEN "110011000000" => table_out <= 3983;
			WHEN "110011000001" => table_out <= 3983;
			WHEN "110011000010" => table_out <= 3983;
			WHEN "110011000011" => table_out <= 3983;
			WHEN "110011000100" => table_out <= 3983;
			WHEN "110011000101" => table_out <= 3984;
			WHEN "110011000110" => table_out <= 3984;
			WHEN "110011000111" => table_out <= 3984;
			WHEN "110011001000" => table_out <= 3984;
			WHEN "110011001001" => table_out <= 3984;
			WHEN "110011001010" => table_out <= 3984;
			WHEN "110011001011" => table_out <= 3985;
			WHEN "110011001100" => table_out <= 3985;
			WHEN "110011001101" => table_out <= 3985;
			WHEN "110011001110" => table_out <= 3985;
			WHEN "110011001111" => table_out <= 3985;
			WHEN "110011010000" => table_out <= 3985;
			WHEN "110011010001" => table_out <= 3985;
			WHEN "110011010010" => table_out <= 3986;
			WHEN "110011010011" => table_out <= 3986;
			WHEN "110011010100" => table_out <= 3986;
			WHEN "110011010101" => table_out <= 3986;
			WHEN "110011010110" => table_out <= 3986;
			WHEN "110011010111" => table_out <= 3986;
			WHEN "110011011000" => table_out <= 3986;
			WHEN "110011011001" => table_out <= 3987;
			WHEN "110011011010" => table_out <= 3987;
			WHEN "110011011011" => table_out <= 3987;
			WHEN "110011011100" => table_out <= 3987;
			WHEN "110011011101" => table_out <= 3987;
			WHEN "110011011110" => table_out <= 3987;
			WHEN "110011011111" => table_out <= 3988;
			WHEN "110011100000" => table_out <= 3988;
			WHEN "110011100001" => table_out <= 3988;
			WHEN "110011100010" => table_out <= 3988;
			WHEN "110011100011" => table_out <= 3988;
			WHEN "110011100100" => table_out <= 3988;
			WHEN "110011100101" => table_out <= 3988;
			WHEN "110011100110" => table_out <= 3989;
			WHEN "110011100111" => table_out <= 3989;
			WHEN "110011101000" => table_out <= 3989;
			WHEN "110011101001" => table_out <= 3989;
			WHEN "110011101010" => table_out <= 3989;
			WHEN "110011101011" => table_out <= 3989;
			WHEN "110011101100" => table_out <= 3989;
			WHEN "110011101101" => table_out <= 3990;
			WHEN "110011101110" => table_out <= 3990;
			WHEN "110011101111" => table_out <= 3990;
			WHEN "110011110000" => table_out <= 3990;
			WHEN "110011110001" => table_out <= 3990;
			WHEN "110011110010" => table_out <= 3990;
			WHEN "110011110011" => table_out <= 3990;
			WHEN "110011110100" => table_out <= 3991;
			WHEN "110011110101" => table_out <= 3991;
			WHEN "110011110110" => table_out <= 3991;
			WHEN "110011110111" => table_out <= 3991;
			WHEN "110011111000" => table_out <= 3991;
			WHEN "110011111001" => table_out <= 3991;
			WHEN "110011111010" => table_out <= 3992;
			WHEN "110011111011" => table_out <= 3992;
			WHEN "110011111100" => table_out <= 3992;
			WHEN "110011111101" => table_out <= 3992;
			WHEN "110011111110" => table_out <= 3992;
			WHEN "110011111111" => table_out <= 3992;
			WHEN "110100000000" => table_out <= 3992;
			WHEN "110100000001" => table_out <= 3993;
			WHEN "110100000010" => table_out <= 3993;
			WHEN "110100000011" => table_out <= 3993;
			WHEN "110100000100" => table_out <= 3993;
			WHEN "110100000101" => table_out <= 3993;
			WHEN "110100000110" => table_out <= 3993;
			WHEN "110100000111" => table_out <= 3993;
			WHEN "110100001000" => table_out <= 3994;
			WHEN "110100001001" => table_out <= 3994;
			WHEN "110100001010" => table_out <= 3994;
			WHEN "110100001011" => table_out <= 3994;
			WHEN "110100001100" => table_out <= 3994;
			WHEN "110100001101" => table_out <= 3994;
			WHEN "110100001110" => table_out <= 3994;
			WHEN "110100001111" => table_out <= 3995;
			WHEN "110100010000" => table_out <= 3995;
			WHEN "110100010001" => table_out <= 3995;
			WHEN "110100010010" => table_out <= 3995;
			WHEN "110100010011" => table_out <= 3995;
			WHEN "110100010100" => table_out <= 3995;
			WHEN "110100010101" => table_out <= 3996;
			WHEN "110100010110" => table_out <= 3996;
			WHEN "110100010111" => table_out <= 3996;
			WHEN "110100011000" => table_out <= 3996;
			WHEN "110100011001" => table_out <= 3996;
			WHEN "110100011010" => table_out <= 3996;
			WHEN "110100011011" => table_out <= 3996;
			WHEN "110100011100" => table_out <= 3997;
			WHEN "110100011101" => table_out <= 3997;
			WHEN "110100011110" => table_out <= 3997;
			WHEN "110100011111" => table_out <= 3997;
			WHEN "110100100000" => table_out <= 3997;
			WHEN "110100100001" => table_out <= 3997;
			WHEN "110100100010" => table_out <= 3997;
			WHEN "110100100011" => table_out <= 3998;
			WHEN "110100100100" => table_out <= 3998;
			WHEN "110100100101" => table_out <= 3998;
			WHEN "110100100110" => table_out <= 3998;
			WHEN "110100100111" => table_out <= 3998;
			WHEN "110100101000" => table_out <= 3998;
			WHEN "110100101001" => table_out <= 3998;
			WHEN "110100101010" => table_out <= 3999;
			WHEN "110100101011" => table_out <= 3999;
			WHEN "110100101100" => table_out <= 3999;
			WHEN "110100101101" => table_out <= 3999;
			WHEN "110100101110" => table_out <= 3999;
			WHEN "110100101111" => table_out <= 3999;
			WHEN "110100110000" => table_out <= 3999;
			WHEN "110100110001" => table_out <= 4000;
			WHEN "110100110010" => table_out <= 4000;
			WHEN "110100110011" => table_out <= 4000;
			WHEN "110100110100" => table_out <= 4000;
			WHEN "110100110101" => table_out <= 4000;
			WHEN "110100110110" => table_out <= 4000;
			WHEN "110100110111" => table_out <= 4000;
			WHEN "110100111000" => table_out <= 4001;
			WHEN "110100111001" => table_out <= 4001;
			WHEN "110100111010" => table_out <= 4001;
			WHEN "110100111011" => table_out <= 4001;
			WHEN "110100111100" => table_out <= 4001;
			WHEN "110100111101" => table_out <= 4001;
			WHEN "110100111110" => table_out <= 4002;
			WHEN "110100111111" => table_out <= 4002;
			WHEN "110101000000" => table_out <= 4002;
			WHEN "110101000001" => table_out <= 4002;
			WHEN "110101000010" => table_out <= 4002;
			WHEN "110101000011" => table_out <= 4002;
			WHEN "110101000100" => table_out <= 4002;
			WHEN "110101000101" => table_out <= 4003;
			WHEN "110101000110" => table_out <= 4003;
			WHEN "110101000111" => table_out <= 4003;
			WHEN "110101001000" => table_out <= 4003;
			WHEN "110101001001" => table_out <= 4003;
			WHEN "110101001010" => table_out <= 4003;
			WHEN "110101001011" => table_out <= 4003;
			WHEN "110101001100" => table_out <= 4004;
			WHEN "110101001101" => table_out <= 4004;
			WHEN "110101001110" => table_out <= 4004;
			WHEN "110101001111" => table_out <= 4004;
			WHEN "110101010000" => table_out <= 4004;
			WHEN "110101010001" => table_out <= 4004;
			WHEN "110101010010" => table_out <= 4004;
			WHEN "110101010011" => table_out <= 4005;
			WHEN "110101010100" => table_out <= 4005;
			WHEN "110101010101" => table_out <= 4005;
			WHEN "110101010110" => table_out <= 4005;
			WHEN "110101010111" => table_out <= 4005;
			WHEN "110101011000" => table_out <= 4005;
			WHEN "110101011001" => table_out <= 4005;
			WHEN "110101011010" => table_out <= 4006;
			WHEN "110101011011" => table_out <= 4006;
			WHEN "110101011100" => table_out <= 4006;
			WHEN "110101011101" => table_out <= 4006;
			WHEN "110101011110" => table_out <= 4006;
			WHEN "110101011111" => table_out <= 4006;
			WHEN "110101100000" => table_out <= 4006;
			WHEN "110101100001" => table_out <= 4007;
			WHEN "110101100010" => table_out <= 4007;
			WHEN "110101100011" => table_out <= 4007;
			WHEN "110101100100" => table_out <= 4007;
			WHEN "110101100101" => table_out <= 4007;
			WHEN "110101100110" => table_out <= 4007;
			WHEN "110101100111" => table_out <= 4007;
			WHEN "110101101000" => table_out <= 4008;
			WHEN "110101101001" => table_out <= 4008;
			WHEN "110101101010" => table_out <= 4008;
			WHEN "110101101011" => table_out <= 4008;
			WHEN "110101101100" => table_out <= 4008;
			WHEN "110101101101" => table_out <= 4008;
			WHEN "110101101110" => table_out <= 4008;
			WHEN "110101101111" => table_out <= 4009;
			WHEN "110101110000" => table_out <= 4009;
			WHEN "110101110001" => table_out <= 4009;
			WHEN "110101110010" => table_out <= 4009;
			WHEN "110101110011" => table_out <= 4009;
			WHEN "110101110100" => table_out <= 4009;
			WHEN "110101110101" => table_out <= 4009;
			WHEN "110101110110" => table_out <= 4010;
			WHEN "110101110111" => table_out <= 4010;
			WHEN "110101111000" => table_out <= 4010;
			WHEN "110101111001" => table_out <= 4010;
			WHEN "110101111010" => table_out <= 4010;
			WHEN "110101111011" => table_out <= 4010;
			WHEN "110101111100" => table_out <= 4010;
			WHEN "110101111101" => table_out <= 4011;
			WHEN "110101111110" => table_out <= 4011;
			WHEN "110101111111" => table_out <= 4011;
			WHEN "110110000000" => table_out <= 4011;
			WHEN "110110000001" => table_out <= 4011;
			WHEN "110110000010" => table_out <= 4011;
			WHEN "110110000011" => table_out <= 4011;
			WHEN "110110000100" => table_out <= 4012;
			WHEN "110110000101" => table_out <= 4012;
			WHEN "110110000110" => table_out <= 4012;
			WHEN "110110000111" => table_out <= 4012;
			WHEN "110110001000" => table_out <= 4012;
			WHEN "110110001001" => table_out <= 4012;
			WHEN "110110001010" => table_out <= 4012;
			WHEN "110110001011" => table_out <= 4013;
			WHEN "110110001100" => table_out <= 4013;
			WHEN "110110001101" => table_out <= 4013;
			WHEN "110110001110" => table_out <= 4013;
			WHEN "110110001111" => table_out <= 4013;
			WHEN "110110010000" => table_out <= 4013;
			WHEN "110110010001" => table_out <= 4013;
			WHEN "110110010010" => table_out <= 4014;
			WHEN "110110010011" => table_out <= 4014;
			WHEN "110110010100" => table_out <= 4014;
			WHEN "110110010101" => table_out <= 4014;
			WHEN "110110010110" => table_out <= 4014;
			WHEN "110110010111" => table_out <= 4014;
			WHEN "110110011000" => table_out <= 4014;
			WHEN "110110011001" => table_out <= 4015;
			WHEN "110110011010" => table_out <= 4015;
			WHEN "110110011011" => table_out <= 4015;
			WHEN "110110011100" => table_out <= 4015;
			WHEN "110110011101" => table_out <= 4015;
			WHEN "110110011110" => table_out <= 4015;
			WHEN "110110011111" => table_out <= 4015;
			WHEN "110110100000" => table_out <= 4016;
			WHEN "110110100001" => table_out <= 4016;
			WHEN "110110100010" => table_out <= 4016;
			WHEN "110110100011" => table_out <= 4016;
			WHEN "110110100100" => table_out <= 4016;
			WHEN "110110100101" => table_out <= 4016;
			WHEN "110110100110" => table_out <= 4016;
			WHEN "110110100111" => table_out <= 4017;
			WHEN "110110101000" => table_out <= 4017;
			WHEN "110110101001" => table_out <= 4017;
			WHEN "110110101010" => table_out <= 4017;
			WHEN "110110101011" => table_out <= 4017;
			WHEN "110110101100" => table_out <= 4017;
			WHEN "110110101101" => table_out <= 4017;
			WHEN "110110101110" => table_out <= 4018;
			WHEN "110110101111" => table_out <= 4018;
			WHEN "110110110000" => table_out <= 4018;
			WHEN "110110110001" => table_out <= 4018;
			WHEN "110110110010" => table_out <= 4018;
			WHEN "110110110011" => table_out <= 4018;
			WHEN "110110110100" => table_out <= 4018;
			WHEN "110110110101" => table_out <= 4018;
			WHEN "110110110110" => table_out <= 4019;
			WHEN "110110110111" => table_out <= 4019;
			WHEN "110110111000" => table_out <= 4019;
			WHEN "110110111001" => table_out <= 4019;
			WHEN "110110111010" => table_out <= 4019;
			WHEN "110110111011" => table_out <= 4019;
			WHEN "110110111100" => table_out <= 4019;
			WHEN "110110111101" => table_out <= 4020;
			WHEN "110110111110" => table_out <= 4020;
			WHEN "110110111111" => table_out <= 4020;
			WHEN "110111000000" => table_out <= 4020;
			WHEN "110111000001" => table_out <= 4020;
			WHEN "110111000010" => table_out <= 4020;
			WHEN "110111000011" => table_out <= 4020;
			WHEN "110111000100" => table_out <= 4021;
			WHEN "110111000101" => table_out <= 4021;
			WHEN "110111000110" => table_out <= 4021;
			WHEN "110111000111" => table_out <= 4021;
			WHEN "110111001000" => table_out <= 4021;
			WHEN "110111001001" => table_out <= 4021;
			WHEN "110111001010" => table_out <= 4021;
			WHEN "110111001011" => table_out <= 4022;
			WHEN "110111001100" => table_out <= 4022;
			WHEN "110111001101" => table_out <= 4022;
			WHEN "110111001110" => table_out <= 4022;
			WHEN "110111001111" => table_out <= 4022;
			WHEN "110111010000" => table_out <= 4022;
			WHEN "110111010001" => table_out <= 4022;
			WHEN "110111010010" => table_out <= 4023;
			WHEN "110111010011" => table_out <= 4023;
			WHEN "110111010100" => table_out <= 4023;
			WHEN "110111010101" => table_out <= 4023;
			WHEN "110111010110" => table_out <= 4023;
			WHEN "110111010111" => table_out <= 4023;
			WHEN "110111011000" => table_out <= 4023;
			WHEN "110111011001" => table_out <= 4024;
			WHEN "110111011010" => table_out <= 4024;
			WHEN "110111011011" => table_out <= 4024;
			WHEN "110111011100" => table_out <= 4024;
			WHEN "110111011101" => table_out <= 4024;
			WHEN "110111011110" => table_out <= 4024;
			WHEN "110111011111" => table_out <= 4024;
			WHEN "110111100000" => table_out <= 4024;
			WHEN "110111100001" => table_out <= 4025;
			WHEN "110111100010" => table_out <= 4025;
			WHEN "110111100011" => table_out <= 4025;
			WHEN "110111100100" => table_out <= 4025;
			WHEN "110111100101" => table_out <= 4025;
			WHEN "110111100110" => table_out <= 4025;
			WHEN "110111100111" => table_out <= 4025;
			WHEN "110111101000" => table_out <= 4026;
			WHEN "110111101001" => table_out <= 4026;
			WHEN "110111101010" => table_out <= 4026;
			WHEN "110111101011" => table_out <= 4026;
			WHEN "110111101100" => table_out <= 4026;
			WHEN "110111101101" => table_out <= 4026;
			WHEN "110111101110" => table_out <= 4026;
			WHEN "110111101111" => table_out <= 4027;
			WHEN "110111110000" => table_out <= 4027;
			WHEN "110111110001" => table_out <= 4027;
			WHEN "110111110010" => table_out <= 4027;
			WHEN "110111110011" => table_out <= 4027;
			WHEN "110111110100" => table_out <= 4027;
			WHEN "110111110101" => table_out <= 4027;
			WHEN "110111110110" => table_out <= 4028;
			WHEN "110111110111" => table_out <= 4028;
			WHEN "110111111000" => table_out <= 4028;
			WHEN "110111111001" => table_out <= 4028;
			WHEN "110111111010" => table_out <= 4028;
			WHEN "110111111011" => table_out <= 4028;
			WHEN "110111111100" => table_out <= 4028;
			WHEN "110111111101" => table_out <= 4028;
			WHEN "110111111110" => table_out <= 4029;
			WHEN "110111111111" => table_out <= 4029;
			WHEN "111000000000" => table_out <= 4029;
			WHEN "111000000001" => table_out <= 4029;
			WHEN "111000000010" => table_out <= 4029;
			WHEN "111000000011" => table_out <= 4029;
			WHEN "111000000100" => table_out <= 4029;
			WHEN "111000000101" => table_out <= 4030;
			WHEN "111000000110" => table_out <= 4030;
			WHEN "111000000111" => table_out <= 4030;
			WHEN "111000001000" => table_out <= 4030;
			WHEN "111000001001" => table_out <= 4030;
			WHEN "111000001010" => table_out <= 4030;
			WHEN "111000001011" => table_out <= 4030;
			WHEN "111000001100" => table_out <= 4031;
			WHEN "111000001101" => table_out <= 4031;
			WHEN "111000001110" => table_out <= 4031;
			WHEN "111000001111" => table_out <= 4031;
			WHEN "111000010000" => table_out <= 4031;
			WHEN "111000010001" => table_out <= 4031;
			WHEN "111000010010" => table_out <= 4031;
			WHEN "111000010011" => table_out <= 4031;
			WHEN "111000010100" => table_out <= 4032;
			WHEN "111000010101" => table_out <= 4032;
			WHEN "111000010110" => table_out <= 4032;
			WHEN "111000010111" => table_out <= 4032;
			WHEN "111000011000" => table_out <= 4032;
			WHEN "111000011001" => table_out <= 4032;
			WHEN "111000011010" => table_out <= 4032;
			WHEN "111000011011" => table_out <= 4033;
			WHEN "111000011100" => table_out <= 4033;
			WHEN "111000011101" => table_out <= 4033;
			WHEN "111000011110" => table_out <= 4033;
			WHEN "111000011111" => table_out <= 4033;
			WHEN "111000100000" => table_out <= 4033;
			WHEN "111000100001" => table_out <= 4033;
			WHEN "111000100010" => table_out <= 4034;
			WHEN "111000100011" => table_out <= 4034;
			WHEN "111000100100" => table_out <= 4034;
			WHEN "111000100101" => table_out <= 4034;
			WHEN "111000100110" => table_out <= 4034;
			WHEN "111000100111" => table_out <= 4034;
			WHEN "111000101000" => table_out <= 4034;
			WHEN "111000101001" => table_out <= 4034;
			WHEN "111000101010" => table_out <= 4035;
			WHEN "111000101011" => table_out <= 4035;
			WHEN "111000101100" => table_out <= 4035;
			WHEN "111000101101" => table_out <= 4035;
			WHEN "111000101110" => table_out <= 4035;
			WHEN "111000101111" => table_out <= 4035;
			WHEN "111000110000" => table_out <= 4035;
			WHEN "111000110001" => table_out <= 4036;
			WHEN "111000110010" => table_out <= 4036;
			WHEN "111000110011" => table_out <= 4036;
			WHEN "111000110100" => table_out <= 4036;
			WHEN "111000110101" => table_out <= 4036;
			WHEN "111000110110" => table_out <= 4036;
			WHEN "111000110111" => table_out <= 4036;
			WHEN "111000111000" => table_out <= 4037;
			WHEN "111000111001" => table_out <= 4037;
			WHEN "111000111010" => table_out <= 4037;
			WHEN "111000111011" => table_out <= 4037;
			WHEN "111000111100" => table_out <= 4037;
			WHEN "111000111101" => table_out <= 4037;
			WHEN "111000111110" => table_out <= 4037;
			WHEN "111000111111" => table_out <= 4037;
			WHEN "111001000000" => table_out <= 4038;
			WHEN "111001000001" => table_out <= 4038;
			WHEN "111001000010" => table_out <= 4038;
			WHEN "111001000011" => table_out <= 4038;
			WHEN "111001000100" => table_out <= 4038;
			WHEN "111001000101" => table_out <= 4038;
			WHEN "111001000110" => table_out <= 4038;
			WHEN "111001000111" => table_out <= 4039;
			WHEN "111001001000" => table_out <= 4039;
			WHEN "111001001001" => table_out <= 4039;
			WHEN "111001001010" => table_out <= 4039;
			WHEN "111001001011" => table_out <= 4039;
			WHEN "111001001100" => table_out <= 4039;
			WHEN "111001001101" => table_out <= 4039;
			WHEN "111001001110" => table_out <= 4039;
			WHEN "111001001111" => table_out <= 4040;
			WHEN "111001010000" => table_out <= 4040;
			WHEN "111001010001" => table_out <= 4040;
			WHEN "111001010010" => table_out <= 4040;
			WHEN "111001010011" => table_out <= 4040;
			WHEN "111001010100" => table_out <= 4040;
			WHEN "111001010101" => table_out <= 4040;
			WHEN "111001010110" => table_out <= 4041;
			WHEN "111001010111" => table_out <= 4041;
			WHEN "111001011000" => table_out <= 4041;
			WHEN "111001011001" => table_out <= 4041;
			WHEN "111001011010" => table_out <= 4041;
			WHEN "111001011011" => table_out <= 4041;
			WHEN "111001011100" => table_out <= 4041;
			WHEN "111001011101" => table_out <= 4042;
			WHEN "111001011110" => table_out <= 4042;
			WHEN "111001011111" => table_out <= 4042;
			WHEN "111001100000" => table_out <= 4042;
			WHEN "111001100001" => table_out <= 4042;
			WHEN "111001100010" => table_out <= 4042;
			WHEN "111001100011" => table_out <= 4042;
			WHEN "111001100100" => table_out <= 4042;
			WHEN "111001100101" => table_out <= 4043;
			WHEN "111001100110" => table_out <= 4043;
			WHEN "111001100111" => table_out <= 4043;
			WHEN "111001101000" => table_out <= 4043;
			WHEN "111001101001" => table_out <= 4043;
			WHEN "111001101010" => table_out <= 4043;
			WHEN "111001101011" => table_out <= 4043;
			WHEN "111001101100" => table_out <= 4044;
			WHEN "111001101101" => table_out <= 4044;
			WHEN "111001101110" => table_out <= 4044;
			WHEN "111001101111" => table_out <= 4044;
			WHEN "111001110000" => table_out <= 4044;
			WHEN "111001110001" => table_out <= 4044;
			WHEN "111001110010" => table_out <= 4044;
			WHEN "111001110011" => table_out <= 4044;
			WHEN "111001110100" => table_out <= 4045;
			WHEN "111001110101" => table_out <= 4045;
			WHEN "111001110110" => table_out <= 4045;
			WHEN "111001110111" => table_out <= 4045;
			WHEN "111001111000" => table_out <= 4045;
			WHEN "111001111001" => table_out <= 4045;
			WHEN "111001111010" => table_out <= 4045;
			WHEN "111001111011" => table_out <= 4046;
			WHEN "111001111100" => table_out <= 4046;
			WHEN "111001111101" => table_out <= 4046;
			WHEN "111001111110" => table_out <= 4046;
			WHEN "111001111111" => table_out <= 4046;
			WHEN "111010000000" => table_out <= 4046;
			WHEN "111010000001" => table_out <= 4046;
			WHEN "111010000010" => table_out <= 4046;
			WHEN "111010000011" => table_out <= 4047;
			WHEN "111010000100" => table_out <= 4047;
			WHEN "111010000101" => table_out <= 4047;
			WHEN "111010000110" => table_out <= 4047;
			WHEN "111010000111" => table_out <= 4047;
			WHEN "111010001000" => table_out <= 4047;
			WHEN "111010001001" => table_out <= 4047;
			WHEN "111010001010" => table_out <= 4047;
			WHEN "111010001011" => table_out <= 4048;
			WHEN "111010001100" => table_out <= 4048;
			WHEN "111010001101" => table_out <= 4048;
			WHEN "111010001110" => table_out <= 4048;
			WHEN "111010001111" => table_out <= 4048;
			WHEN "111010010000" => table_out <= 4048;
			WHEN "111010010001" => table_out <= 4048;
			WHEN "111010010010" => table_out <= 4049;
			WHEN "111010010011" => table_out <= 4049;
			WHEN "111010010100" => table_out <= 4049;
			WHEN "111010010101" => table_out <= 4049;
			WHEN "111010010110" => table_out <= 4049;
			WHEN "111010010111" => table_out <= 4049;
			WHEN "111010011000" => table_out <= 4049;
			WHEN "111010011001" => table_out <= 4049;
			WHEN "111010011010" => table_out <= 4050;
			WHEN "111010011011" => table_out <= 4050;
			WHEN "111010011100" => table_out <= 4050;
			WHEN "111010011101" => table_out <= 4050;
			WHEN "111010011110" => table_out <= 4050;
			WHEN "111010011111" => table_out <= 4050;
			WHEN "111010100000" => table_out <= 4050;
			WHEN "111010100001" => table_out <= 4051;
			WHEN "111010100010" => table_out <= 4051;
			WHEN "111010100011" => table_out <= 4051;
			WHEN "111010100100" => table_out <= 4051;
			WHEN "111010100101" => table_out <= 4051;
			WHEN "111010100110" => table_out <= 4051;
			WHEN "111010100111" => table_out <= 4051;
			WHEN "111010101000" => table_out <= 4051;
			WHEN "111010101001" => table_out <= 4052;
			WHEN "111010101010" => table_out <= 4052;
			WHEN "111010101011" => table_out <= 4052;
			WHEN "111010101100" => table_out <= 4052;
			WHEN "111010101101" => table_out <= 4052;
			WHEN "111010101110" => table_out <= 4052;
			WHEN "111010101111" => table_out <= 4052;
			WHEN "111010110000" => table_out <= 4052;
			WHEN "111010110001" => table_out <= 4053;
			WHEN "111010110010" => table_out <= 4053;
			WHEN "111010110011" => table_out <= 4053;
			WHEN "111010110100" => table_out <= 4053;
			WHEN "111010110101" => table_out <= 4053;
			WHEN "111010110110" => table_out <= 4053;
			WHEN "111010110111" => table_out <= 4053;
			WHEN "111010111000" => table_out <= 4054;
			WHEN "111010111001" => table_out <= 4054;
			WHEN "111010111010" => table_out <= 4054;
			WHEN "111010111011" => table_out <= 4054;
			WHEN "111010111100" => table_out <= 4054;
			WHEN "111010111101" => table_out <= 4054;
			WHEN "111010111110" => table_out <= 4054;
			WHEN "111010111111" => table_out <= 4054;
			WHEN "111011000000" => table_out <= 4055;
			WHEN "111011000001" => table_out <= 4055;
			WHEN "111011000010" => table_out <= 4055;
			WHEN "111011000011" => table_out <= 4055;
			WHEN "111011000100" => table_out <= 4055;
			WHEN "111011000101" => table_out <= 4055;
			WHEN "111011000110" => table_out <= 4055;
			WHEN "111011000111" => table_out <= 4055;
			WHEN "111011001000" => table_out <= 4056;
			WHEN "111011001001" => table_out <= 4056;
			WHEN "111011001010" => table_out <= 4056;
			WHEN "111011001011" => table_out <= 4056;
			WHEN "111011001100" => table_out <= 4056;
			WHEN "111011001101" => table_out <= 4056;
			WHEN "111011001110" => table_out <= 4056;
			WHEN "111011001111" => table_out <= 4057;
			WHEN "111011010000" => table_out <= 4057;
			WHEN "111011010001" => table_out <= 4057;
			WHEN "111011010010" => table_out <= 4057;
			WHEN "111011010011" => table_out <= 4057;
			WHEN "111011010100" => table_out <= 4057;
			WHEN "111011010101" => table_out <= 4057;
			WHEN "111011010110" => table_out <= 4057;
			WHEN "111011010111" => table_out <= 4058;
			WHEN "111011011000" => table_out <= 4058;
			WHEN "111011011001" => table_out <= 4058;
			WHEN "111011011010" => table_out <= 4058;
			WHEN "111011011011" => table_out <= 4058;
			WHEN "111011011100" => table_out <= 4058;
			WHEN "111011011101" => table_out <= 4058;
			WHEN "111011011110" => table_out <= 4058;
			WHEN "111011011111" => table_out <= 4059;
			WHEN "111011100000" => table_out <= 4059;
			WHEN "111011100001" => table_out <= 4059;
			WHEN "111011100010" => table_out <= 4059;
			WHEN "111011100011" => table_out <= 4059;
			WHEN "111011100100" => table_out <= 4059;
			WHEN "111011100101" => table_out <= 4059;
			WHEN "111011100110" => table_out <= 4060;
			WHEN "111011100111" => table_out <= 4060;
			WHEN "111011101000" => table_out <= 4060;
			WHEN "111011101001" => table_out <= 4060;
			WHEN "111011101010" => table_out <= 4060;
			WHEN "111011101011" => table_out <= 4060;
			WHEN "111011101100" => table_out <= 4060;
			WHEN "111011101101" => table_out <= 4060;
			WHEN "111011101110" => table_out <= 4061;
			WHEN "111011101111" => table_out <= 4061;
			WHEN "111011110000" => table_out <= 4061;
			WHEN "111011110001" => table_out <= 4061;
			WHEN "111011110010" => table_out <= 4061;
			WHEN "111011110011" => table_out <= 4061;
			WHEN "111011110100" => table_out <= 4061;
			WHEN "111011110101" => table_out <= 4061;
			WHEN "111011110110" => table_out <= 4062;
			WHEN "111011110111" => table_out <= 4062;
			WHEN "111011111000" => table_out <= 4062;
			WHEN "111011111001" => table_out <= 4062;
			WHEN "111011111010" => table_out <= 4062;
			WHEN "111011111011" => table_out <= 4062;
			WHEN "111011111100" => table_out <= 4062;
			WHEN "111011111101" => table_out <= 4062;
			WHEN "111011111110" => table_out <= 4063;
			WHEN "111011111111" => table_out <= 4063;
			WHEN "111100000000" => table_out <= 4063;
			WHEN "111100000001" => table_out <= 4063;
			WHEN "111100000010" => table_out <= 4063;
			WHEN "111100000011" => table_out <= 4063;
			WHEN "111100000100" => table_out <= 4063;
			WHEN "111100000101" => table_out <= 4063;
			WHEN "111100000110" => table_out <= 4064;
			WHEN "111100000111" => table_out <= 4064;
			WHEN "111100001000" => table_out <= 4064;
			WHEN "111100001001" => table_out <= 4064;
			WHEN "111100001010" => table_out <= 4064;
			WHEN "111100001011" => table_out <= 4064;
			WHEN "111100001100" => table_out <= 4064;
			WHEN "111100001101" => table_out <= 4065;
			WHEN "111100001110" => table_out <= 4065;
			WHEN "111100001111" => table_out <= 4065;
			WHEN "111100010000" => table_out <= 4065;
			WHEN "111100010001" => table_out <= 4065;
			WHEN "111100010010" => table_out <= 4065;
			WHEN "111100010011" => table_out <= 4065;
			WHEN "111100010100" => table_out <= 4065;
			WHEN "111100010101" => table_out <= 4066;
			WHEN "111100010110" => table_out <= 4066;
			WHEN "111100010111" => table_out <= 4066;
			WHEN "111100011000" => table_out <= 4066;
			WHEN "111100011001" => table_out <= 4066;
			WHEN "111100011010" => table_out <= 4066;
			WHEN "111100011011" => table_out <= 4066;
			WHEN "111100011100" => table_out <= 4066;
			WHEN "111100011101" => table_out <= 4067;
			WHEN "111100011110" => table_out <= 4067;
			WHEN "111100011111" => table_out <= 4067;
			WHEN "111100100000" => table_out <= 4067;
			WHEN "111100100001" => table_out <= 4067;
			WHEN "111100100010" => table_out <= 4067;
			WHEN "111100100011" => table_out <= 4067;
			WHEN "111100100100" => table_out <= 4067;
			WHEN "111100100101" => table_out <= 4068;
			WHEN "111100100110" => table_out <= 4068;
			WHEN "111100100111" => table_out <= 4068;
			WHEN "111100101000" => table_out <= 4068;
			WHEN "111100101001" => table_out <= 4068;
			WHEN "111100101010" => table_out <= 4068;
			WHEN "111100101011" => table_out <= 4068;
			WHEN "111100101100" => table_out <= 4068;
			WHEN "111100101101" => table_out <= 4069;
			WHEN "111100101110" => table_out <= 4069;
			WHEN "111100101111" => table_out <= 4069;
			WHEN "111100110000" => table_out <= 4069;
			WHEN "111100110001" => table_out <= 4069;
			WHEN "111100110010" => table_out <= 4069;
			WHEN "111100110011" => table_out <= 4069;
			WHEN "111100110100" => table_out <= 4069;
			WHEN "111100110101" => table_out <= 4070;
			WHEN "111100110110" => table_out <= 4070;
			WHEN "111100110111" => table_out <= 4070;
			WHEN "111100111000" => table_out <= 4070;
			WHEN "111100111001" => table_out <= 4070;
			WHEN "111100111010" => table_out <= 4070;
			WHEN "111100111011" => table_out <= 4070;
			WHEN "111100111100" => table_out <= 4070;
			WHEN "111100111101" => table_out <= 4071;
			WHEN "111100111110" => table_out <= 4071;
			WHEN "111100111111" => table_out <= 4071;
			WHEN "111101000000" => table_out <= 4071;
			WHEN "111101000001" => table_out <= 4071;
			WHEN "111101000010" => table_out <= 4071;
			WHEN "111101000011" => table_out <= 4071;
			WHEN "111101000100" => table_out <= 4071;
			WHEN "111101000101" => table_out <= 4072;
			WHEN "111101000110" => table_out <= 4072;
			WHEN "111101000111" => table_out <= 4072;
			WHEN "111101001000" => table_out <= 4072;
			WHEN "111101001001" => table_out <= 4072;
			WHEN "111101001010" => table_out <= 4072;
			WHEN "111101001011" => table_out <= 4072;
			WHEN "111101001100" => table_out <= 4073;
			WHEN "111101001101" => table_out <= 4073;
			WHEN "111101001110" => table_out <= 4073;
			WHEN "111101001111" => table_out <= 4073;
			WHEN "111101010000" => table_out <= 4073;
			WHEN "111101010001" => table_out <= 4073;
			WHEN "111101010010" => table_out <= 4073;
			WHEN "111101010011" => table_out <= 4073;
			WHEN "111101010100" => table_out <= 4074;
			WHEN "111101010101" => table_out <= 4074;
			WHEN "111101010110" => table_out <= 4074;
			WHEN "111101010111" => table_out <= 4074;
			WHEN "111101011000" => table_out <= 4074;
			WHEN "111101011001" => table_out <= 4074;
			WHEN "111101011010" => table_out <= 4074;
			WHEN "111101011011" => table_out <= 4074;
			WHEN "111101011100" => table_out <= 4075;
			WHEN "111101011101" => table_out <= 4075;
			WHEN "111101011110" => table_out <= 4075;
			WHEN "111101011111" => table_out <= 4075;
			WHEN "111101100000" => table_out <= 4075;
			WHEN "111101100001" => table_out <= 4075;
			WHEN "111101100010" => table_out <= 4075;
			WHEN "111101100011" => table_out <= 4075;
			WHEN "111101100100" => table_out <= 4076;
			WHEN "111101100101" => table_out <= 4076;
			WHEN "111101100110" => table_out <= 4076;
			WHEN "111101100111" => table_out <= 4076;
			WHEN "111101101000" => table_out <= 4076;
			WHEN "111101101001" => table_out <= 4076;
			WHEN "111101101010" => table_out <= 4076;
			WHEN "111101101011" => table_out <= 4076;
			WHEN "111101101100" => table_out <= 4077;
			WHEN "111101101101" => table_out <= 4077;
			WHEN "111101101110" => table_out <= 4077;
			WHEN "111101101111" => table_out <= 4077;
			WHEN "111101110000" => table_out <= 4077;
			WHEN "111101110001" => table_out <= 4077;
			WHEN "111101110010" => table_out <= 4077;
			WHEN "111101110011" => table_out <= 4077;
			WHEN "111101110100" => table_out <= 4078;
			WHEN "111101110101" => table_out <= 4078;
			WHEN "111101110110" => table_out <= 4078;
			WHEN "111101110111" => table_out <= 4078;
			WHEN "111101111000" => table_out <= 4078;
			WHEN "111101111001" => table_out <= 4078;
			WHEN "111101111010" => table_out <= 4078;
			WHEN "111101111011" => table_out <= 4078;
			WHEN "111101111100" => table_out <= 4078;
			WHEN "111101111101" => table_out <= 4079;
			WHEN "111101111110" => table_out <= 4079;
			WHEN "111101111111" => table_out <= 4079;
			WHEN "111110000000" => table_out <= 4079;
			WHEN "111110000001" => table_out <= 4079;
			WHEN "111110000010" => table_out <= 4079;
			WHEN "111110000011" => table_out <= 4079;
			WHEN "111110000100" => table_out <= 4079;
			WHEN "111110000101" => table_out <= 4080;
			WHEN "111110000110" => table_out <= 4080;
			WHEN "111110000111" => table_out <= 4080;
			WHEN "111110001000" => table_out <= 4080;
			WHEN "111110001001" => table_out <= 4080;
			WHEN "111110001010" => table_out <= 4080;
			WHEN "111110001011" => table_out <= 4080;
			WHEN "111110001100" => table_out <= 4080;
			WHEN "111110001101" => table_out <= 4081;
			WHEN "111110001110" => table_out <= 4081;
			WHEN "111110001111" => table_out <= 4081;
			WHEN "111110010000" => table_out <= 4081;
			WHEN "111110010001" => table_out <= 4081;
			WHEN "111110010010" => table_out <= 4081;
			WHEN "111110010011" => table_out <= 4081;
			WHEN "111110010100" => table_out <= 4081;
			WHEN "111110010101" => table_out <= 4082;
			WHEN "111110010110" => table_out <= 4082;
			WHEN "111110010111" => table_out <= 4082;
			WHEN "111110011000" => table_out <= 4082;
			WHEN "111110011001" => table_out <= 4082;
			WHEN "111110011010" => table_out <= 4082;
			WHEN "111110011011" => table_out <= 4082;
			WHEN "111110011100" => table_out <= 4082;
			WHEN "111110011101" => table_out <= 4083;
			WHEN "111110011110" => table_out <= 4083;
			WHEN "111110011111" => table_out <= 4083;
			WHEN "111110100000" => table_out <= 4083;
			WHEN "111110100001" => table_out <= 4083;
			WHEN "111110100010" => table_out <= 4083;
			WHEN "111110100011" => table_out <= 4083;
			WHEN "111110100100" => table_out <= 4083;
			WHEN "111110100101" => table_out <= 4084;
			WHEN "111110100110" => table_out <= 4084;
			WHEN "111110100111" => table_out <= 4084;
			WHEN "111110101000" => table_out <= 4084;
			WHEN "111110101001" => table_out <= 4084;
			WHEN "111110101010" => table_out <= 4084;
			WHEN "111110101011" => table_out <= 4084;
			WHEN "111110101100" => table_out <= 4084;
			WHEN "111110101101" => table_out <= 4085;
			WHEN "111110101110" => table_out <= 4085;
			WHEN "111110101111" => table_out <= 4085;
			WHEN "111110110000" => table_out <= 4085;
			WHEN "111110110001" => table_out <= 4085;
			WHEN "111110110010" => table_out <= 4085;
			WHEN "111110110011" => table_out <= 4085;
			WHEN "111110110100" => table_out <= 4085;
			WHEN "111110110101" => table_out <= 4086;
			WHEN "111110110110" => table_out <= 4086;
			WHEN "111110110111" => table_out <= 4086;
			WHEN "111110111000" => table_out <= 4086;
			WHEN "111110111001" => table_out <= 4086;
			WHEN "111110111010" => table_out <= 4086;
			WHEN "111110111011" => table_out <= 4086;
			WHEN "111110111100" => table_out <= 4086;
			WHEN "111110111101" => table_out <= 4087;
			WHEN "111110111110" => table_out <= 4087;
			WHEN "111110111111" => table_out <= 4087;
			WHEN "111111000000" => table_out <= 4087;
			WHEN "111111000001" => table_out <= 4087;
			WHEN "111111000010" => table_out <= 4087;
			WHEN "111111000011" => table_out <= 4087;
			WHEN "111111000100" => table_out <= 4087;
			WHEN "111111000101" => table_out <= 4087;
			WHEN "111111000110" => table_out <= 4088;
			WHEN "111111000111" => table_out <= 4088;
			WHEN "111111001000" => table_out <= 4088;
			WHEN "111111001001" => table_out <= 4088;
			WHEN "111111001010" => table_out <= 4088;
			WHEN "111111001011" => table_out <= 4088;
			WHEN "111111001100" => table_out <= 4088;
			WHEN "111111001101" => table_out <= 4088;
			WHEN "111111001110" => table_out <= 4089;
			WHEN "111111001111" => table_out <= 4089;
			WHEN "111111010000" => table_out <= 4089;
			WHEN "111111010001" => table_out <= 4089;
			WHEN "111111010010" => table_out <= 4089;
			WHEN "111111010011" => table_out <= 4089;
			WHEN "111111010100" => table_out <= 4089;
			WHEN "111111010101" => table_out <= 4089;
			WHEN "111111010110" => table_out <= 4090;
			WHEN "111111010111" => table_out <= 4090;
			WHEN "111111011000" => table_out <= 4090;
			WHEN "111111011001" => table_out <= 4090;
			WHEN "111111011010" => table_out <= 4090;
			WHEN "111111011011" => table_out <= 4090;
			WHEN "111111011100" => table_out <= 4090;
			WHEN "111111011101" => table_out <= 4090;
			WHEN "111111011110" => table_out <= 4091;
			WHEN "111111011111" => table_out <= 4091;
			WHEN "111111100000" => table_out <= 4091;
			WHEN "111111100001" => table_out <= 4091;
			WHEN "111111100010" => table_out <= 4091;
			WHEN "111111100011" => table_out <= 4091;
			WHEN "111111100100" => table_out <= 4091;
			WHEN "111111100101" => table_out <= 4091;
			WHEN "111111100110" => table_out <= 4091;
			WHEN "111111100111" => table_out <= 4092;
			WHEN "111111101000" => table_out <= 4092;
			WHEN "111111101001" => table_out <= 4092;
			WHEN "111111101010" => table_out <= 4092;
			WHEN "111111101011" => table_out <= 4092;
			WHEN "111111101100" => table_out <= 4092;
			WHEN "111111101101" => table_out <= 4092;
			WHEN "111111101110" => table_out <= 4092;
			WHEN "111111101111" => table_out <= 4093;
			WHEN "111111110000" => table_out <= 4093;
			WHEN "111111110001" => table_out <= 4093;
			WHEN "111111110010" => table_out <= 4093;
			WHEN "111111110011" => table_out <= 4093;
			WHEN "111111110100" => table_out <= 4093;
			WHEN "111111110101" => table_out <= 4093;
			WHEN "111111110110" => table_out <= 4093;
			WHEN "111111110111" => table_out <= 4094;
			WHEN "111111111000" => table_out <= 4094;
			WHEN "111111111001" => table_out <= 4094;
			WHEN "111111111010" => table_out <= 4094;
			WHEN "111111111011" => table_out <= 4094;
			WHEN "111111111100" => table_out <= 4094;
			WHEN "111111111101" => table_out <= 4094;
			WHEN "111111111110" => table_out <= 4094;
			WHEN "111111111111" => table_out <= 4095;
			WHEN OTHERS => table_out <= 0;
		END CASE;
	END PROCESS;
END Behavior;